library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity compteur_led is
  port(
    sysclk        :in  std_logic;
    sw            :in  std_logic_vector(3 downto 0);
    btn           :in  std_logic_vector(3 downto 0);
    led           :out std_logic_vector(3 downto 0)
  );
end compteur_led;

architecture behaviour of compteur_led is
  signal counter : unsigned(31 downto 0) := to_unsigned(0, 32); 
  
component PS7
  port (
     DMA0DATYPE : out std_logic_vector(1 downto 0);
     DMA0DAVALID : out std_ulogic;
     DMA0DRREADY : out std_ulogic;
     DMA0RSTN : out std_ulogic;
     DMA1DATYPE : out std_logic_vector(1 downto 0);
     DMA1DAVALID : out std_ulogic;
     DMA1DRREADY : out std_ulogic;
     DMA1RSTN : out std_ulogic;
     DMA2DATYPE : out std_logic_vector(1 downto 0);
     DMA2DAVALID : out std_ulogic;
     DMA2DRREADY : out std_ulogic;
     DMA2RSTN : out std_ulogic;
     DMA3DATYPE : out std_logic_vector(1 downto 0);
     DMA3DAVALID : out std_ulogic;
     DMA3DRREADY : out std_ulogic;
     DMA3RSTN : out std_ulogic;
     EMIOCAN0PHYTX : out std_ulogic;
     EMIOCAN1PHYTX : out std_ulogic;
     EMIOENET0GMIITXD : out std_logic_vector(7 downto 0);
     EMIOENET0GMIITXEN : out std_ulogic;
     EMIOENET0GMIITXER : out std_ulogic;
     EMIOENET0MDIOMDC : out std_ulogic;
     EMIOENET0MDIOO : out std_ulogic;
     EMIOENET0MDIOTN : out std_ulogic;
     EMIOENET0PTPDELAYREQRX : out std_ulogic;
     EMIOENET0PTPDELAYREQTX : out std_ulogic;
     EMIOENET0PTPPDELAYREQRX : out std_ulogic;
     EMIOENET0PTPPDELAYREQTX : out std_ulogic;
     EMIOENET0PTPPDELAYRESPRX : out std_ulogic;
     EMIOENET0PTPPDELAYRESPTX : out std_ulogic;
     EMIOENET0PTPSYNCFRAMERX : out std_ulogic;
     EMIOENET0PTPSYNCFRAMETX : out std_ulogic;
     EMIOENET0SOFRX : out std_ulogic;
     EMIOENET0SOFTX : out std_ulogic;
     EMIOENET1GMIITXD : out std_logic_vector(7 downto 0);
     EMIOENET1GMIITXEN : out std_ulogic;
     EMIOENET1GMIITXER : out std_ulogic;
     EMIOENET1MDIOMDC : out std_ulogic;
     EMIOENET1MDIOO : out std_ulogic;
     EMIOENET1MDIOTN : out std_ulogic;
     EMIOENET1PTPDELAYREQRX : out std_ulogic;
     EMIOENET1PTPDELAYREQTX : out std_ulogic;
     EMIOENET1PTPPDELAYREQRX : out std_ulogic;
     EMIOENET1PTPPDELAYREQTX : out std_ulogic;
     EMIOENET1PTPPDELAYRESPRX : out std_ulogic;
     EMIOENET1PTPPDELAYRESPTX : out std_ulogic;
     EMIOENET1PTPSYNCFRAMERX : out std_ulogic;
     EMIOENET1PTPSYNCFRAMETX : out std_ulogic;
     EMIOENET1SOFRX : out std_ulogic;
     EMIOENET1SOFTX : out std_ulogic;
     EMIOGPIOO : out std_logic_vector(63 downto 0);
     EMIOGPIOTN : out std_logic_vector(63 downto 0);
     EMIOI2C0SCLO : out std_ulogic;
     EMIOI2C0SCLTN : out std_ulogic;
     EMIOI2C0SDAO : out std_ulogic;
     EMIOI2C0SDATN : out std_ulogic;
     EMIOI2C1SCLO : out std_ulogic;
     EMIOI2C1SCLTN : out std_ulogic;
     EMIOI2C1SDAO : out std_ulogic;
     EMIOI2C1SDATN : out std_ulogic;
     EMIOPJTAGTDO : out std_ulogic;
     EMIOPJTAGTDTN : out std_ulogic;
     EMIOSDIO0BUSPOW : out std_ulogic;
     EMIOSDIO0BUSVOLT : out std_logic_vector(2 downto 0);
     EMIOSDIO0CLK : out std_ulogic;
     EMIOSDIO0CMDO : out std_ulogic;
     EMIOSDIO0CMDTN : out std_ulogic;
     EMIOSDIO0DATAO : out std_logic_vector(3 downto 0);
     EMIOSDIO0DATATN : out std_logic_vector(3 downto 0);
     EMIOSDIO0LED : out std_ulogic;
     EMIOSDIO1BUSPOW : out std_ulogic;
     EMIOSDIO1BUSVOLT : out std_logic_vector(2 downto 0);
     EMIOSDIO1CLK : out std_ulogic;
     EMIOSDIO1CMDO : out std_ulogic;
     EMIOSDIO1CMDTN : out std_ulogic;
     EMIOSDIO1DATAO : out std_logic_vector(3 downto 0);
     EMIOSDIO1DATATN : out std_logic_vector(3 downto 0);
     EMIOSDIO1LED : out std_ulogic;
     EMIOSPI0MO : out std_ulogic;
     EMIOSPI0MOTN : out std_ulogic;
     EMIOSPI0SCLKO : out std_ulogic;
     EMIOSPI0SCLKTN : out std_ulogic;
     EMIOSPI0SO : out std_ulogic;
     EMIOSPI0SSNTN : out std_ulogic;
     EMIOSPI0SSON : out std_logic_vector(2 downto 0);
     EMIOSPI0STN : out std_ulogic;
     EMIOSPI1MO : out std_ulogic;
     EMIOSPI1MOTN : out std_ulogic;
     EMIOSPI1SCLKO : out std_ulogic;
     EMIOSPI1SCLKTN : out std_ulogic;
     EMIOSPI1SO : out std_ulogic;
     EMIOSPI1SSNTN : out std_ulogic;
     EMIOSPI1SSON : out std_logic_vector(2 downto 0);
     EMIOSPI1STN : out std_ulogic;
     EMIOTRACECTL : out std_ulogic;
     EMIOTRACEDATA : out std_logic_vector(31 downto 0);
     EMIOTTC0WAVEO : out std_logic_vector(2 downto 0);
     EMIOTTC1WAVEO : out std_logic_vector(2 downto 0);
     EMIOUART0DTRN : out std_ulogic;
     EMIOUART0RTSN : out std_ulogic;
     EMIOUART0TX : out std_ulogic;
     EMIOUART1DTRN : out std_ulogic;
     EMIOUART1RTSN : out std_ulogic;
     EMIOUART1TX : out std_ulogic;
     EMIOUSB0PORTINDCTL : out std_logic_vector(1 downto 0);
     EMIOUSB0VBUSPWRSELECT : out std_ulogic;
     EMIOUSB1PORTINDCTL : out std_logic_vector(1 downto 0);
     EMIOUSB1VBUSPWRSELECT : out std_ulogic;
     EMIOWDTRSTO : out std_ulogic;
     EVENTEVENTO : out std_ulogic;
     EVENTSTANDBYWFE : out std_logic_vector(1 downto 0);
     EVENTSTANDBYWFI : out std_logic_vector(1 downto 0);
     FCLKCLK : out std_logic_vector(3 downto 0);
     FCLKRESETN : out std_logic_vector(3 downto 0);
     FTMTF2PTRIGACK : out std_logic_vector(3 downto 0);
     FTMTP2FDEBUG : out std_logic_vector(31 downto 0);
     FTMTP2FTRIG : out std_logic_vector(3 downto 0);
     IRQP2F : out std_logic_vector(28 downto 0);
     MAXIGP0ARADDR : out std_logic_vector(31 downto 0);
     MAXIGP0ARBURST : out std_logic_vector(1 downto 0);
     MAXIGP0ARCACHE : out std_logic_vector(3 downto 0);
     MAXIGP0ARESETN : out std_ulogic;
     MAXIGP0ARID : out std_logic_vector(11 downto 0);
     MAXIGP0ARLEN : out std_logic_vector(3 downto 0);
     MAXIGP0ARLOCK : out std_logic_vector(1 downto 0);
     MAXIGP0ARPROT : out std_logic_vector(2 downto 0);
     MAXIGP0ARQOS : out std_logic_vector(3 downto 0);
     MAXIGP0ARSIZE : out std_logic_vector(1 downto 0);
     MAXIGP0ARVALID : out std_ulogic;
     MAXIGP0AWADDR : out std_logic_vector(31 downto 0);
     MAXIGP0AWBURST : out std_logic_vector(1 downto 0);
     MAXIGP0AWCACHE : out std_logic_vector(3 downto 0);
     MAXIGP0AWID : out std_logic_vector(11 downto 0);
     MAXIGP0AWLEN : out std_logic_vector(3 downto 0);
     MAXIGP0AWLOCK : out std_logic_vector(1 downto 0);
     MAXIGP0AWPROT : out std_logic_vector(2 downto 0);
     MAXIGP0AWQOS : out std_logic_vector(3 downto 0);
     MAXIGP0AWSIZE : out std_logic_vector(1 downto 0);
     MAXIGP0AWVALID : out std_ulogic;
     MAXIGP0BREADY : out std_ulogic;
     MAXIGP0RREADY : out std_ulogic;
     MAXIGP0WDATA : out std_logic_vector(31 downto 0);
     MAXIGP0WID : out std_logic_vector(11 downto 0);
     MAXIGP0WLAST : out std_ulogic;
     MAXIGP0WSTRB : out std_logic_vector(3 downto 0);
     MAXIGP0WVALID : out std_ulogic;
     MAXIGP1ARADDR : out std_logic_vector(31 downto 0);
     MAXIGP1ARBURST : out std_logic_vector(1 downto 0);
     MAXIGP1ARCACHE : out std_logic_vector(3 downto 0);
     MAXIGP1ARESETN : out std_ulogic;
     MAXIGP1ARID : out std_logic_vector(11 downto 0);
     MAXIGP1ARLEN : out std_logic_vector(3 downto 0);
     MAXIGP1ARLOCK : out std_logic_vector(1 downto 0);
     MAXIGP1ARPROT : out std_logic_vector(2 downto 0);
     MAXIGP1ARQOS : out std_logic_vector(3 downto 0);
     MAXIGP1ARSIZE : out std_logic_vector(1 downto 0);
     MAXIGP1ARVALID : out std_ulogic;
     MAXIGP1AWADDR : out std_logic_vector(31 downto 0);
     MAXIGP1AWBURST : out std_logic_vector(1 downto 0);
     MAXIGP1AWCACHE : out std_logic_vector(3 downto 0);
     MAXIGP1AWID : out std_logic_vector(11 downto 0);
     MAXIGP1AWLEN : out std_logic_vector(3 downto 0);
     MAXIGP1AWLOCK : out std_logic_vector(1 downto 0);
     MAXIGP1AWPROT : out std_logic_vector(2 downto 0);
     MAXIGP1AWQOS : out std_logic_vector(3 downto 0);
     MAXIGP1AWSIZE : out std_logic_vector(1 downto 0);
     MAXIGP1AWVALID : out std_ulogic;
     MAXIGP1BREADY : out std_ulogic;
     MAXIGP1RREADY : out std_ulogic;
     MAXIGP1WDATA : out std_logic_vector(31 downto 0);
     MAXIGP1WID : out std_logic_vector(11 downto 0);
     MAXIGP1WLAST : out std_ulogic;
     MAXIGP1WSTRB : out std_logic_vector(3 downto 0);
     MAXIGP1WVALID : out std_ulogic;
     SAXIACPARESETN : out std_ulogic;
     SAXIACPARREADY : out std_ulogic;
     SAXIACPAWREADY : out std_ulogic;
     SAXIACPBID : out std_logic_vector(2 downto 0);
     SAXIACPBRESP : out std_logic_vector(1 downto 0);
     SAXIACPBVALID : out std_ulogic;
     SAXIACPRDATA : out std_logic_vector(63 downto 0);
     SAXIACPRID : out std_logic_vector(2 downto 0);
     SAXIACPRLAST : out std_ulogic;
     SAXIACPRRESP : out std_logic_vector(1 downto 0);
     SAXIACPRVALID : out std_ulogic;
     SAXIACPWREADY : out std_ulogic;
     SAXIGP0ARESETN : out std_ulogic;
     SAXIGP0ARREADY : out std_ulogic;
     SAXIGP0AWREADY : out std_ulogic;
     SAXIGP0BID : out std_logic_vector(5 downto 0);
     SAXIGP0BRESP : out std_logic_vector(1 downto 0);
     SAXIGP0BVALID : out std_ulogic;
     SAXIGP0RDATA : out std_logic_vector(31 downto 0);
     SAXIGP0RID : out std_logic_vector(5 downto 0);
     SAXIGP0RLAST : out std_ulogic;
     SAXIGP0RRESP : out std_logic_vector(1 downto 0);
     SAXIGP0RVALID : out std_ulogic;
     SAXIGP0WREADY : out std_ulogic;
     SAXIGP1ARESETN : out std_ulogic;
     SAXIGP1ARREADY : out std_ulogic;
     SAXIGP1AWREADY : out std_ulogic;
     SAXIGP1BID : out std_logic_vector(5 downto 0);
     SAXIGP1BRESP : out std_logic_vector(1 downto 0);
     SAXIGP1BVALID : out std_ulogic;
     SAXIGP1RDATA : out std_logic_vector(31 downto 0);
     SAXIGP1RID : out std_logic_vector(5 downto 0);
     SAXIGP1RLAST : out std_ulogic;
     SAXIGP1RRESP : out std_logic_vector(1 downto 0);
     SAXIGP1RVALID : out std_ulogic;
     SAXIGP1WREADY : out std_ulogic;
     SAXIHP0ARESETN : out std_ulogic;
     SAXIHP0ARREADY : out std_ulogic;
     SAXIHP0AWREADY : out std_ulogic;
     SAXIHP0BID : out std_logic_vector(5 downto 0);
     SAXIHP0BRESP : out std_logic_vector(1 downto 0);
     SAXIHP0BVALID : out std_ulogic;
     SAXIHP0RACOUNT : out std_logic_vector(2 downto 0);
     SAXIHP0RCOUNT : out std_logic_vector(7 downto 0);
     SAXIHP0RDATA : out std_logic_vector(63 downto 0);
     SAXIHP0RID : out std_logic_vector(5 downto 0);
     SAXIHP0RLAST : out std_ulogic;
     SAXIHP0RRESP : out std_logic_vector(1 downto 0);
     SAXIHP0RVALID : out std_ulogic;
     SAXIHP0WACOUNT : out std_logic_vector(5 downto 0);
     SAXIHP0WCOUNT : out std_logic_vector(7 downto 0);
     SAXIHP0WREADY : out std_ulogic;
     SAXIHP1ARESETN : out std_ulogic;
     SAXIHP1ARREADY : out std_ulogic;
     SAXIHP1AWREADY : out std_ulogic;
     SAXIHP1BID : out std_logic_vector(5 downto 0);
     SAXIHP1BRESP : out std_logic_vector(1 downto 0);
     SAXIHP1BVALID : out std_ulogic;
     SAXIHP1RACOUNT : out std_logic_vector(2 downto 0);
     SAXIHP1RCOUNT : out std_logic_vector(7 downto 0);
     SAXIHP1RDATA : out std_logic_vector(63 downto 0);
     SAXIHP1RID : out std_logic_vector(5 downto 0);
     SAXIHP1RLAST : out std_ulogic;
     SAXIHP1RRESP : out std_logic_vector(1 downto 0);
     SAXIHP1RVALID : out std_ulogic;
     SAXIHP1WACOUNT : out std_logic_vector(5 downto 0);
     SAXIHP1WCOUNT : out std_logic_vector(7 downto 0);
     SAXIHP1WREADY : out std_ulogic;
     SAXIHP2ARESETN : out std_ulogic;
     SAXIHP2ARREADY : out std_ulogic;
     SAXIHP2AWREADY : out std_ulogic;
     SAXIHP2BID : out std_logic_vector(5 downto 0);
     SAXIHP2BRESP : out std_logic_vector(1 downto 0);
     SAXIHP2BVALID : out std_ulogic;
     SAXIHP2RACOUNT : out std_logic_vector(2 downto 0);
     SAXIHP2RCOUNT : out std_logic_vector(7 downto 0);
     SAXIHP2RDATA : out std_logic_vector(63 downto 0);
     SAXIHP2RID : out std_logic_vector(5 downto 0);
     SAXIHP2RLAST : out std_ulogic;
     SAXIHP2RRESP : out std_logic_vector(1 downto 0);
     SAXIHP2RVALID : out std_ulogic;
     SAXIHP2WACOUNT : out std_logic_vector(5 downto 0);
     SAXIHP2WCOUNT : out std_logic_vector(7 downto 0);
     SAXIHP2WREADY : out std_ulogic;
     SAXIHP3ARESETN : out std_ulogic;
     SAXIHP3ARREADY : out std_ulogic;
     SAXIHP3AWREADY : out std_ulogic;
     SAXIHP3BID : out std_logic_vector(5 downto 0);
     SAXIHP3BRESP : out std_logic_vector(1 downto 0);
     SAXIHP3BVALID : out std_ulogic;
     SAXIHP3RACOUNT : out std_logic_vector(2 downto 0);
     SAXIHP3RCOUNT : out std_logic_vector(7 downto 0);
     SAXIHP3RDATA : out std_logic_vector(63 downto 0);
     SAXIHP3RID : out std_logic_vector(5 downto 0);
     SAXIHP3RLAST : out std_ulogic;
     SAXIHP3RRESP : out std_logic_vector(1 downto 0);
     SAXIHP3RVALID : out std_ulogic;
     SAXIHP3WACOUNT : out std_logic_vector(5 downto 0);
     SAXIHP3WCOUNT : out std_logic_vector(7 downto 0);
     SAXIHP3WREADY : out std_ulogic;
     DDRA : inout std_logic_vector(14 downto 0);
     DDRBA : inout std_logic_vector(2 downto 0);
     DDRCASB : inout std_ulogic;
     DDRCKE : inout std_ulogic;
     DDRCKN : inout std_ulogic;
     DDRCKP : inout std_ulogic;
     DDRCSB : inout std_ulogic;
     DDRDM : inout std_logic_vector(3 downto 0);
     DDRDQ : inout std_logic_vector(31 downto 0);
     DDRDQSN : inout std_logic_vector(3 downto 0);
     DDRDQSP : inout std_logic_vector(3 downto 0);
     DDRDRSTB : inout std_ulogic;
     DDRODT : inout std_ulogic;
     DDRRASB : inout std_ulogic;
     DDRVRN : inout std_ulogic;
     DDRVRP : inout std_ulogic;
     DDRWEB : inout std_ulogic;
     MIO : inout std_logic_vector(53 downto 0);
     PSCLK : inout std_ulogic;
     PSPORB : inout std_ulogic;
     PSSRSTB : inout std_ulogic;
     DDRARB : in std_logic_vector(3 downto 0);
     DMA0ACLK : in std_ulogic;
     DMA0DAREADY : in std_ulogic;
     DMA0DRLAST : in std_ulogic;
     DMA0DRTYPE : in std_logic_vector(1 downto 0);
     DMA0DRVALID : in std_ulogic;
     DMA1ACLK : in std_ulogic;
     DMA1DAREADY : in std_ulogic;
     DMA1DRLAST : in std_ulogic;
     DMA1DRTYPE : in std_logic_vector(1 downto 0);
     DMA1DRVALID : in std_ulogic;
     DMA2ACLK : in std_ulogic;
     DMA2DAREADY : in std_ulogic;
     DMA2DRLAST : in std_ulogic;
     DMA2DRTYPE : in std_logic_vector(1 downto 0);
     DMA2DRVALID : in std_ulogic;
     DMA3ACLK : in std_ulogic;
     DMA3DAREADY : in std_ulogic;
     DMA3DRLAST : in std_ulogic;
     DMA3DRTYPE : in std_logic_vector(1 downto 0);
     DMA3DRVALID : in std_ulogic;
     EMIOCAN0PHYRX : in std_ulogic;
     EMIOCAN1PHYRX : in std_ulogic;
     EMIOENET0EXTINTIN : in std_ulogic;
     EMIOENET0GMIICOL : in std_ulogic;
     EMIOENET0GMIICRS : in std_ulogic;
     EMIOENET0GMIIRXCLK : in std_ulogic;
     EMIOENET0GMIIRXD : in std_logic_vector(7 downto 0);
     EMIOENET0GMIIRXDV : in std_ulogic;
     EMIOENET0GMIIRXER : in std_ulogic;
     EMIOENET0GMIITXCLK : in std_ulogic;
     EMIOENET0MDIOI : in std_ulogic;
     EMIOENET1EXTINTIN : in std_ulogic;
     EMIOENET1GMIICOL : in std_ulogic;
     EMIOENET1GMIICRS : in std_ulogic;
     EMIOENET1GMIIRXCLK : in std_ulogic;
     EMIOENET1GMIIRXD : in std_logic_vector(7 downto 0);
     EMIOENET1GMIIRXDV : in std_ulogic;
     EMIOENET1GMIIRXER : in std_ulogic;
     EMIOENET1GMIITXCLK : in std_ulogic;
     EMIOENET1MDIOI : in std_ulogic;
     EMIOGPIOI : in std_logic_vector(63 downto 0);
     EMIOI2C0SCLI : in std_ulogic;
     EMIOI2C0SDAI : in std_ulogic;
     EMIOI2C1SCLI : in std_ulogic;
     EMIOI2C1SDAI : in std_ulogic;
     EMIOPJTAGTCK : in std_ulogic;
     EMIOPJTAGTDI : in std_ulogic;
     EMIOPJTAGTMS : in std_ulogic;
     EMIOSDIO0CDN : in std_ulogic;
     EMIOSDIO0CLKFB : in std_ulogic;
     EMIOSDIO0CMDI : in std_ulogic;
     EMIOSDIO0DATAI : in std_logic_vector(3 downto 0);
     EMIOSDIO0WP : in std_ulogic;
     EMIOSDIO1CDN : in std_ulogic;
     EMIOSDIO1CLKFB : in std_ulogic;
     EMIOSDIO1CMDI : in std_ulogic;
     EMIOSDIO1DATAI : in std_logic_vector(3 downto 0);
     EMIOSDIO1WP : in std_ulogic;
     EMIOSPI0MI : in std_ulogic;
     EMIOSPI0SCLKI : in std_ulogic;
     EMIOSPI0SI : in std_ulogic;
     EMIOSPI0SSIN : in std_ulogic;
     EMIOSPI1MI : in std_ulogic;
     EMIOSPI1SCLKI : in std_ulogic;
     EMIOSPI1SI : in std_ulogic;
     EMIOSPI1SSIN : in std_ulogic;
     EMIOSRAMINTIN : in std_ulogic;
     EMIOTRACECLK : in std_ulogic;
     EMIOTTC0CLKI : in std_logic_vector(2 downto 0);
     EMIOTTC1CLKI : in std_logic_vector(2 downto 0);
     EMIOUART0CTSN : in std_ulogic;
     EMIOUART0DCDN : in std_ulogic;
     EMIOUART0DSRN : in std_ulogic;
     EMIOUART0RIN : in std_ulogic;
     EMIOUART0RX : in std_ulogic;
     EMIOUART1CTSN : in std_ulogic;
     EMIOUART1DCDN : in std_ulogic;
     EMIOUART1DSRN : in std_ulogic;
     EMIOUART1RIN : in std_ulogic;
     EMIOUART1RX : in std_ulogic;
     EMIOUSB0VBUSPWRFAULT : in std_ulogic;
     EMIOUSB1VBUSPWRFAULT : in std_ulogic;
     EMIOWDTCLKI : in std_ulogic;
     EVENTEVENTI : in std_ulogic;
     FCLKCLKTRIGN : in std_logic_vector(3 downto 0);
     FPGAIDLEN : in std_ulogic;
     FTMDTRACEINATID : in std_logic_vector(3 downto 0);
     FTMDTRACEINCLOCK : in std_ulogic;
     FTMDTRACEINDATA : in std_logic_vector(31 downto 0);
     FTMDTRACEINVALID : in std_ulogic;
     FTMTF2PDEBUG : in std_logic_vector(31 downto 0);
     FTMTF2PTRIG : in std_logic_vector(3 downto 0);
     FTMTP2FTRIGACK : in std_logic_vector(3 downto 0);
     IRQF2P : in std_logic_vector(19 downto 0);
     MAXIGP0ACLK : in std_ulogic;
     MAXIGP0ARREADY : in std_ulogic;
     MAXIGP0AWREADY : in std_ulogic;
     MAXIGP0BID : in std_logic_vector(11 downto 0);
     MAXIGP0BRESP : in std_logic_vector(1 downto 0);
     MAXIGP0BVALID : in std_ulogic;
     MAXIGP0RDATA : in std_logic_vector(31 downto 0);
     MAXIGP0RID : in std_logic_vector(11 downto 0);
     MAXIGP0RLAST : in std_ulogic;
     MAXIGP0RRESP : in std_logic_vector(1 downto 0);
     MAXIGP0RVALID : in std_ulogic;
     MAXIGP0WREADY : in std_ulogic;
     MAXIGP1ACLK : in std_ulogic;
     MAXIGP1ARREADY : in std_ulogic;
     MAXIGP1AWREADY : in std_ulogic;
     MAXIGP1BID : in std_logic_vector(11 downto 0);
     MAXIGP1BRESP : in std_logic_vector(1 downto 0);
     MAXIGP1BVALID : in std_ulogic;
     MAXIGP1RDATA : in std_logic_vector(31 downto 0);
     MAXIGP1RID : in std_logic_vector(11 downto 0);
     MAXIGP1RLAST : in std_ulogic;
     MAXIGP1RRESP : in std_logic_vector(1 downto 0);
     MAXIGP1RVALID : in std_ulogic;
     MAXIGP1WREADY : in std_ulogic;
     SAXIACPACLK : in std_ulogic;
     SAXIACPARADDR : in std_logic_vector(31 downto 0);
     SAXIACPARBURST : in std_logic_vector(1 downto 0);
     SAXIACPARCACHE : in std_logic_vector(3 downto 0);
     SAXIACPARID : in std_logic_vector(2 downto 0);
     SAXIACPARLEN : in std_logic_vector(3 downto 0);
     SAXIACPARLOCK : in std_logic_vector(1 downto 0);
     SAXIACPARPROT : in std_logic_vector(2 downto 0);
     SAXIACPARQOS : in std_logic_vector(3 downto 0);
     SAXIACPARSIZE : in std_logic_vector(1 downto 0);
     SAXIACPARUSER : in std_logic_vector(4 downto 0);
     SAXIACPARVALID : in std_ulogic;
     SAXIACPAWADDR : in std_logic_vector(31 downto 0);
     SAXIACPAWBURST : in std_logic_vector(1 downto 0);
     SAXIACPAWCACHE : in std_logic_vector(3 downto 0);
     SAXIACPAWID : in std_logic_vector(2 downto 0);
     SAXIACPAWLEN : in std_logic_vector(3 downto 0);
     SAXIACPAWLOCK : in std_logic_vector(1 downto 0);
     SAXIACPAWPROT : in std_logic_vector(2 downto 0);
     SAXIACPAWQOS : in std_logic_vector(3 downto 0);
     SAXIACPAWSIZE : in std_logic_vector(1 downto 0);
     SAXIACPAWUSER : in std_logic_vector(4 downto 0);
     SAXIACPAWVALID : in std_ulogic;
     SAXIACPBREADY : in std_ulogic;
     SAXIACPRREADY : in std_ulogic;
     SAXIACPWDATA : in std_logic_vector(63 downto 0);
     SAXIACPWID : in std_logic_vector(2 downto 0);
     SAXIACPWLAST : in std_ulogic;
     SAXIACPWSTRB : in std_logic_vector(7 downto 0);
     SAXIACPWVALID : in std_ulogic;
     SAXIGP0ACLK : in std_ulogic;
     SAXIGP0ARADDR : in std_logic_vector(31 downto 0);
     SAXIGP0ARBURST : in std_logic_vector(1 downto 0);
     SAXIGP0ARCACHE : in std_logic_vector(3 downto 0);
     SAXIGP0ARID : in std_logic_vector(5 downto 0);
     SAXIGP0ARLEN : in std_logic_vector(3 downto 0);
     SAXIGP0ARLOCK : in std_logic_vector(1 downto 0);
     SAXIGP0ARPROT : in std_logic_vector(2 downto 0);
     SAXIGP0ARQOS : in std_logic_vector(3 downto 0);
     SAXIGP0ARSIZE : in std_logic_vector(1 downto 0);
     SAXIGP0ARVALID : in std_ulogic;
     SAXIGP0AWADDR : in std_logic_vector(31 downto 0);
     SAXIGP0AWBURST : in std_logic_vector(1 downto 0);
     SAXIGP0AWCACHE : in std_logic_vector(3 downto 0);
     SAXIGP0AWID : in std_logic_vector(5 downto 0);
     SAXIGP0AWLEN : in std_logic_vector(3 downto 0);
     SAXIGP0AWLOCK : in std_logic_vector(1 downto 0);
     SAXIGP0AWPROT : in std_logic_vector(2 downto 0);
     SAXIGP0AWQOS : in std_logic_vector(3 downto 0);
     SAXIGP0AWSIZE : in std_logic_vector(1 downto 0);
     SAXIGP0AWVALID : in std_ulogic;
     SAXIGP0BREADY : in std_ulogic;
     SAXIGP0RREADY : in std_ulogic;
     SAXIGP0WDATA : in std_logic_vector(31 downto 0);
     SAXIGP0WID : in std_logic_vector(5 downto 0);
     SAXIGP0WLAST : in std_ulogic;
     SAXIGP0WSTRB : in std_logic_vector(3 downto 0);
     SAXIGP0WVALID : in std_ulogic;
     SAXIGP1ACLK : in std_ulogic;
     SAXIGP1ARADDR : in std_logic_vector(31 downto 0);
     SAXIGP1ARBURST : in std_logic_vector(1 downto 0);
     SAXIGP1ARCACHE : in std_logic_vector(3 downto 0);
     SAXIGP1ARID : in std_logic_vector(5 downto 0);
     SAXIGP1ARLEN : in std_logic_vector(3 downto 0);
     SAXIGP1ARLOCK : in std_logic_vector(1 downto 0);
     SAXIGP1ARPROT : in std_logic_vector(2 downto 0);
     SAXIGP1ARQOS : in std_logic_vector(3 downto 0);
     SAXIGP1ARSIZE : in std_logic_vector(1 downto 0);
     SAXIGP1ARVALID : in std_ulogic;
     SAXIGP1AWADDR : in std_logic_vector(31 downto 0);
     SAXIGP1AWBURST : in std_logic_vector(1 downto 0);
     SAXIGP1AWCACHE : in std_logic_vector(3 downto 0);
     SAXIGP1AWID : in std_logic_vector(5 downto 0);
     SAXIGP1AWLEN : in std_logic_vector(3 downto 0);
     SAXIGP1AWLOCK : in std_logic_vector(1 downto 0);
     SAXIGP1AWPROT : in std_logic_vector(2 downto 0);
     SAXIGP1AWQOS : in std_logic_vector(3 downto 0);
     SAXIGP1AWSIZE : in std_logic_vector(1 downto 0);
     SAXIGP1AWVALID : in std_ulogic;
     SAXIGP1BREADY : in std_ulogic;
     SAXIGP1RREADY : in std_ulogic;
     SAXIGP1WDATA : in std_logic_vector(31 downto 0);
     SAXIGP1WID : in std_logic_vector(5 downto 0);
     SAXIGP1WLAST : in std_ulogic;
     SAXIGP1WSTRB : in std_logic_vector(3 downto 0);
     SAXIGP1WVALID : in std_ulogic;
     SAXIHP0ACLK : in std_ulogic;
     SAXIHP0ARADDR : in std_logic_vector(31 downto 0);
     SAXIHP0ARBURST : in std_logic_vector(1 downto 0);
     SAXIHP0ARCACHE : in std_logic_vector(3 downto 0);
     SAXIHP0ARID : in std_logic_vector(5 downto 0);
     SAXIHP0ARLEN : in std_logic_vector(3 downto 0);
     SAXIHP0ARLOCK : in std_logic_vector(1 downto 0);
     SAXIHP0ARPROT : in std_logic_vector(2 downto 0);
     SAXIHP0ARQOS : in std_logic_vector(3 downto 0);
     SAXIHP0ARSIZE : in std_logic_vector(1 downto 0);
     SAXIHP0ARVALID : in std_ulogic;
     SAXIHP0AWADDR : in std_logic_vector(31 downto 0);
     SAXIHP0AWBURST : in std_logic_vector(1 downto 0);
     SAXIHP0AWCACHE : in std_logic_vector(3 downto 0);
     SAXIHP0AWID : in std_logic_vector(5 downto 0);
     SAXIHP0AWLEN : in std_logic_vector(3 downto 0);
     SAXIHP0AWLOCK : in std_logic_vector(1 downto 0);
     SAXIHP0AWPROT : in std_logic_vector(2 downto 0);
     SAXIHP0AWQOS : in std_logic_vector(3 downto 0);
     SAXIHP0AWSIZE : in std_logic_vector(1 downto 0);
     SAXIHP0AWVALID : in std_ulogic;
     SAXIHP0BREADY : in std_ulogic;
     SAXIHP0RDISSUECAP1EN : in std_ulogic;
     SAXIHP0RREADY : in std_ulogic;
     SAXIHP0WDATA : in std_logic_vector(63 downto 0);
     SAXIHP0WID : in std_logic_vector(5 downto 0);
     SAXIHP0WLAST : in std_ulogic;
     SAXIHP0WRISSUECAP1EN : in std_ulogic;
     SAXIHP0WSTRB : in std_logic_vector(7 downto 0);
     SAXIHP0WVALID : in std_ulogic;
     SAXIHP1ACLK : in std_ulogic;
     SAXIHP1ARADDR : in std_logic_vector(31 downto 0);
     SAXIHP1ARBURST : in std_logic_vector(1 downto 0);
     SAXIHP1ARCACHE : in std_logic_vector(3 downto 0);
     SAXIHP1ARID : in std_logic_vector(5 downto 0);
     SAXIHP1ARLEN : in std_logic_vector(3 downto 0);
     SAXIHP1ARLOCK : in std_logic_vector(1 downto 0);
     SAXIHP1ARPROT : in std_logic_vector(2 downto 0);
     SAXIHP1ARQOS : in std_logic_vector(3 downto 0);
     SAXIHP1ARSIZE : in std_logic_vector(1 downto 0);
     SAXIHP1ARVALID : in std_ulogic;
     SAXIHP1AWADDR : in std_logic_vector(31 downto 0);
     SAXIHP1AWBURST : in std_logic_vector(1 downto 0);
     SAXIHP1AWCACHE : in std_logic_vector(3 downto 0);
     SAXIHP1AWID : in std_logic_vector(5 downto 0);
     SAXIHP1AWLEN : in std_logic_vector(3 downto 0);
     SAXIHP1AWLOCK : in std_logic_vector(1 downto 0);
     SAXIHP1AWPROT : in std_logic_vector(2 downto 0);
     SAXIHP1AWQOS : in std_logic_vector(3 downto 0);
     SAXIHP1AWSIZE : in std_logic_vector(1 downto 0);
     SAXIHP1AWVALID : in std_ulogic;
     SAXIHP1BREADY : in std_ulogic;
     SAXIHP1RDISSUECAP1EN : in std_ulogic;
     SAXIHP1RREADY : in std_ulogic;
     SAXIHP1WDATA : in std_logic_vector(63 downto 0);
     SAXIHP1WID : in std_logic_vector(5 downto 0);
     SAXIHP1WLAST : in std_ulogic;
     SAXIHP1WRISSUECAP1EN : in std_ulogic;
     SAXIHP1WSTRB : in std_logic_vector(7 downto 0);
     SAXIHP1WVALID : in std_ulogic;
     SAXIHP2ACLK : in std_ulogic;
     SAXIHP2ARADDR : in std_logic_vector(31 downto 0);
     SAXIHP2ARBURST : in std_logic_vector(1 downto 0);
     SAXIHP2ARCACHE : in std_logic_vector(3 downto 0);
     SAXIHP2ARID : in std_logic_vector(5 downto 0);
     SAXIHP2ARLEN : in std_logic_vector(3 downto 0);
     SAXIHP2ARLOCK : in std_logic_vector(1 downto 0);
     SAXIHP2ARPROT : in std_logic_vector(2 downto 0);
     SAXIHP2ARQOS : in std_logic_vector(3 downto 0);
     SAXIHP2ARSIZE : in std_logic_vector(1 downto 0);
     SAXIHP2ARVALID : in std_ulogic;
     SAXIHP2AWADDR : in std_logic_vector(31 downto 0);
     SAXIHP2AWBURST : in std_logic_vector(1 downto 0);
     SAXIHP2AWCACHE : in std_logic_vector(3 downto 0);
     SAXIHP2AWID : in std_logic_vector(5 downto 0);
     SAXIHP2AWLEN : in std_logic_vector(3 downto 0);
     SAXIHP2AWLOCK : in std_logic_vector(1 downto 0);
     SAXIHP2AWPROT : in std_logic_vector(2 downto 0);
     SAXIHP2AWQOS : in std_logic_vector(3 downto 0);
     SAXIHP2AWSIZE : in std_logic_vector(1 downto 0);
     SAXIHP2AWVALID : in std_ulogic;
     SAXIHP2BREADY : in std_ulogic;
     SAXIHP2RDISSUECAP1EN : in std_ulogic;
     SAXIHP2RREADY : in std_ulogic;
     SAXIHP2WDATA : in std_logic_vector(63 downto 0);
     SAXIHP2WID : in std_logic_vector(5 downto 0);
     SAXIHP2WLAST : in std_ulogic;
     SAXIHP2WRISSUECAP1EN : in std_ulogic;
     SAXIHP2WSTRB : in std_logic_vector(7 downto 0);
     SAXIHP2WVALID : in std_ulogic;
     SAXIHP3ACLK : in std_ulogic;
     SAXIHP3ARADDR : in std_logic_vector(31 downto 0);
     SAXIHP3ARBURST : in std_logic_vector(1 downto 0);
     SAXIHP3ARCACHE : in std_logic_vector(3 downto 0);
     SAXIHP3ARID : in std_logic_vector(5 downto 0);
     SAXIHP3ARLEN : in std_logic_vector(3 downto 0);
     SAXIHP3ARLOCK : in std_logic_vector(1 downto 0);
     SAXIHP3ARPROT : in std_logic_vector(2 downto 0);
     SAXIHP3ARQOS : in std_logic_vector(3 downto 0);
     SAXIHP3ARSIZE : in std_logic_vector(1 downto 0);
     SAXIHP3ARVALID : in std_ulogic;
     SAXIHP3AWADDR : in std_logic_vector(31 downto 0);
     SAXIHP3AWBURST : in std_logic_vector(1 downto 0);
     SAXIHP3AWCACHE : in std_logic_vector(3 downto 0);
     SAXIHP3AWID : in std_logic_vector(5 downto 0);
     SAXIHP3AWLEN : in std_logic_vector(3 downto 0);
     SAXIHP3AWLOCK : in std_logic_vector(1 downto 0);
     SAXIHP3AWPROT : in std_logic_vector(2 downto 0);
     SAXIHP3AWQOS : in std_logic_vector(3 downto 0);
     SAXIHP3AWSIZE : in std_logic_vector(1 downto 0);
     SAXIHP3AWVALID : in std_ulogic;
     SAXIHP3BREADY : in std_ulogic;
     SAXIHP3RDISSUECAP1EN : in std_ulogic;
     SAXIHP3RREADY : in std_ulogic;
     SAXIHP3WDATA : in std_logic_vector(63 downto 0);
     SAXIHP3WID : in std_logic_vector(5 downto 0);
     SAXIHP3WLAST : in std_ulogic;
     SAXIHP3WRISSUECAP1EN : in std_ulogic;
     SAXIHP3WSTRB : in std_logic_vector(7 downto 0);
     SAXIHP3WVALID : in std_ulogic
  );
end component;
--attribute BOX_TYPE of
 -- PS7 : component is "PRIMITIVE";
  
begin
  PS7_inst : PS7
    port map (
	DMA0DATYPE			=> open,		-- out std_logic_vector(1 downto 0);
	DMA0DAVALID			=> open,		-- out std_ulogic;
	DMA0DRREADY			=> open,		-- out std_ulogic;
	DMA0RSTN			=> open,		-- out std_ulogic;
	DMA1DATYPE			=> open,		-- out std_logic_vector(1 downto 0);
	DMA1DAVALID			=> open,		-- out std_ulogic;
	DMA1DRREADY			=> open,		-- out std_ulogic;
	DMA1RSTN			=> open,		-- out std_ulogic;
	DMA2DATYPE			=> open,		-- out std_logic_vector(1 downto 0);
	DMA2DAVALID			=> open,		-- out std_ulogic;
	DMA2DRREADY			=> open,		-- out std_ulogic;
	DMA2RSTN			=> open,		-- out std_ulogic;
	DMA3DATYPE			=> open,		-- out std_logic_vector(1 downto 0);
	DMA3DAVALID			=> open,		-- out std_ulogic;
	DMA3DRREADY			=> open,		-- out std_ulogic;
	DMA3RSTN			=> open,		-- out std_ulogic;
	EMIOCAN0PHYTX			=> open,		-- out std_ulogic;
	EMIOCAN1PHYTX			=> open,		-- out std_ulogic;
	EMIOENET0GMIITXD		=> open,		-- out std_logic_vector(7 downto 0);
	EMIOENET0GMIITXEN		=> open,		-- out std_ulogic;
	EMIOENET0GMIITXER		=> open,		-- out std_ulogic;
	EMIOENET0MDIOMDC		=> open,		-- out std_ulogic;
	EMIOENET0MDIOO			=> open,		-- out std_ulogic;
	EMIOENET0MDIOTN			=> open,		-- out std_ulogic;
	EMIOENET0PTPDELAYREQRX		=> open,		-- out std_ulogic;
	EMIOENET0PTPDELAYREQTX		=> open,		-- out std_ulogic;
	EMIOENET0PTPPDELAYREQRX		=> open,		-- out std_ulogic;
	EMIOENET0PTPPDELAYREQTX		=> open,		-- out std_ulogic;
	EMIOENET0PTPPDELAYRESPRX	=> open,		-- out std_ulogic;
	EMIOENET0PTPPDELAYRESPTX	=> open,		-- out std_ulogic;
	EMIOENET0PTPSYNCFRAMERX		=> open,		-- out std_ulogic;
	EMIOENET0PTPSYNCFRAMETX		=> open,		-- out std_ulogic;
	EMIOENET0SOFRX			=> open,		-- out std_ulogic;
	EMIOENET0SOFTX			=> open,		-- out std_ulogic;
	EMIOENET1GMIITXD		=> open,		-- out std_logic_vector(7 downto 0);
	EMIOENET1GMIITXEN		=> open,		-- out std_ulogic;
	EMIOENET1GMIITXER		=> open,		-- out std_ulogic;
	EMIOENET1MDIOMDC		=> open,		-- out std_ulogic;
	EMIOENET1MDIOO			=> open,		-- out std_ulogic;
	EMIOENET1MDIOTN			=> open,		-- out std_ulogic;
	EMIOENET1PTPDELAYREQRX		=> open,		-- out std_ulogic;
	EMIOENET1PTPDELAYREQTX		=> open,		-- out std_ulogic;
	EMIOENET1PTPPDELAYREQRX		=> open,		-- out std_ulogic;
	EMIOENET1PTPPDELAYREQTX		=> open,		-- out std_ulogic;
	EMIOENET1PTPPDELAYRESPRX	=> open,		-- out std_ulogic;
	EMIOENET1PTPPDELAYRESPTX	=> open,		-- out std_ulogic;
	EMIOENET1PTPSYNCFRAMERX		=> open,		-- out std_ulogic;
	EMIOENET1PTPSYNCFRAMETX		=> open,		-- out std_ulogic;
	EMIOENET1SOFRX			=> open,		-- out std_ulogic;
	EMIOENET1SOFTX			=> open,		-- out std_ulogic;
	EMIOGPIOO			=> open,		-- out std_logic_vector(63 downto 0);
	EMIOGPIOTN			=> open,		-- out std_logic_vector(63 downto 0);
	EMIOI2C0SCLO			=> open,		-- out std_ulogic;
	EMIOI2C0SCLTN			=> open,		-- out std_ulogic;
	EMIOI2C0SDAO			=> open,		-- out std_ulogic;
	EMIOI2C0SDATN			=> open,		-- out std_ulogic;
	EMIOI2C1SCLO			=> open,		-- out std_ulogic;
	EMIOI2C1SCLTN			=> open,		-- out std_ulogic;
	EMIOI2C1SDAO			=> open,		-- out std_ulogic;
	EMIOI2C1SDATN			=> open,		-- out std_ulogic;
	EMIOPJTAGTDO			=> open,		-- out std_ulogic;
	EMIOPJTAGTDTN			=> open,		-- out std_ulogic;
	EMIOSDIO0BUSPOW			=> open,		-- out std_ulogic;
	EMIOSDIO0BUSVOLT		=> open,		-- out std_logic_vector(2 downto 0);
	EMIOSDIO0CLK			=> open,		-- out std_ulogic;
	EMIOSDIO0CMDO			=> open,		-- out std_ulogic;
	EMIOSDIO0CMDTN			=> open,		-- out std_ulogic;
	EMIOSDIO0DATAO			=> open,		-- out std_logic_vector(3 downto 0);
	EMIOSDIO0DATATN			=> open,		-- out std_logic_vector(3 downto 0);
	EMIOSDIO0LED			=> open,		-- out std_ulogic;
	EMIOSDIO1BUSPOW			=> open,		-- out std_ulogic;
	EMIOSDIO1BUSVOLT		=> open,		-- out std_logic_vector(2 downto 0);
	EMIOSDIO1CLK			=> open,		-- out std_ulogic;
	EMIOSDIO1CMDO			=> open,		-- out std_ulogic;
	EMIOSDIO1CMDTN			=> open,		-- out std_ulogic;
	EMIOSDIO1DATAO			=> open,		-- out std_logic_vector(3 downto 0);
	EMIOSDIO1DATATN			=> open,		-- out std_logic_vector(3 downto 0);
	EMIOSDIO1LED			=> open,		-- out std_ulogic;
	EMIOSPI0MO			=> open,		-- out std_ulogic;
	EMIOSPI0MOTN			=> open,		-- out std_ulogic;
	EMIOSPI0SCLKO			=> open,		-- out std_ulogic;
	EMIOSPI0SCLKTN			=> open,		-- out std_ulogic;
	EMIOSPI0SO			=> open,		-- out std_ulogic;
	EMIOSPI0SSNTN			=> open,		-- out std_ulogic;
	EMIOSPI0SSON			=> open,		-- out std_logic_vector(2 downto 0);
	EMIOSPI0STN			=> open,		-- out std_ulogic;
	EMIOSPI1MO			=> open,		-- out std_ulogic;
	EMIOSPI1MOTN			=> open,		-- out std_ulogic;
	EMIOSPI1SCLKO			=> open,		-- out std_ulogic;
	EMIOSPI1SCLKTN			=> open,		-- out std_ulogic;
	EMIOSPI1SO			=> open,		-- out std_ulogic;
	EMIOSPI1SSNTN			=> open,		-- out std_ulogic;
	EMIOSPI1SSON			=> open,		-- out std_logic_vector(2 downto 0);
	EMIOSPI1STN			=> open,		-- out std_ulogic;
	EMIOTRACECTL			=> open,		-- out std_ulogic;
	EMIOTRACEDATA			=> open,		-- out std_logic_vector(31 downto 0);
	EMIOTTC0WAVEO			=> open,		-- out std_logic_vector(2 downto 0);
	EMIOTTC1WAVEO			=> open,		-- out std_logic_vector(2 downto 0);
	EMIOUART0DTRN			=> open,		-- out std_ulogic;
	EMIOUART0RTSN			=> open,		-- out std_ulogic;
	EMIOUART0TX			=> open,		-- out std_ulogic;
	EMIOUART1DTRN			=> open,		-- out std_ulogic;
	EMIOUART1RTSN			=> open,		-- out std_ulogic;
	EMIOUART1TX			=> open,		-- out std_ulogic;
	EMIOUSB0PORTINDCTL		=> open,		-- out std_logic_vector(1 downto 0);
	EMIOUSB0VBUSPWRSELECT		=> open,		-- out std_ulogic;
	EMIOUSB1PORTINDCTL		=> open,		-- out std_logic_vector(1 downto 0);
	EMIOUSB1VBUSPWRSELECT		=> open,		-- out std_ulogic;
	EMIOWDTRSTO			=> open,		-- out std_ulogic;
	EVENTEVENTO			=> open,		-- out std_ulogic;
	EVENTSTANDBYWFE			=> open,		-- out std_logic_vector(1 downto 0);
	EVENTSTANDBYWFI			=> open,		-- out std_logic_vector(1 downto 0);
	FCLKCLK				=> open,		-- out std_logic_vector(3 downto 0);
	FCLKRESETN			=> open,		-- out std_logic_vector(3 downto 0);
	FTMTF2PTRIGACK			=> open,		-- out std_logic_vector(3 downto 0);
	FTMTP2FDEBUG			=> open,		-- out std_logic_vector(31 downto 0);
	FTMTP2FTRIG			=> open,		-- out std_logic_vector(3 downto 0);
	IRQP2F				=> open,		-- out std_logic_vector(28 downto 0);
	MAXIGP0ARADDR			=> open,		-- out std_logic_vector(31 downto 0);
	MAXIGP0ARBURST			=> open,		-- out std_logic_vector(1 downto 0);
	MAXIGP0ARCACHE			=> open,		-- out std_logic_vector(3 downto 0);
	MAXIGP0ARESETN			=> open,		-- out std_ulogic;
	MAXIGP0ARID			=> open,		-- out std_logic_vector(11 downto 0);
	MAXIGP0ARLEN			=> open,		-- out std_logic_vector(3 downto 0);
	MAXIGP0ARLOCK			=> open,		-- out std_logic_vector(1 downto 0);
	MAXIGP0ARPROT			=> open,		-- out std_logic_vector(2 downto 0);
	MAXIGP0ARQOS			=> open,		-- out std_logic_vector(3 downto 0);
	MAXIGP0ARSIZE			=> open,		-- out std_logic_vector(1 downto 0);
	MAXIGP0ARVALID			=> open,		-- out std_ulogic;
	MAXIGP0AWADDR			=> open,		-- out std_logic_vector(31 downto 0);
	MAXIGP0AWBURST			=> open,		-- out std_logic_vector(1 downto 0);
	MAXIGP0AWCACHE			=> open,		-- out std_logic_vector(3 downto 0);
	MAXIGP0AWID			=> open,		-- out std_logic_vector(11 downto 0);
	MAXIGP0AWLEN			=> open,		-- out std_logic_vector(3 downto 0);
	MAXIGP0AWLOCK			=> open,		-- out std_logic_vector(1 downto 0);
	MAXIGP0AWPROT			=> open,		-- out std_logic_vector(2 downto 0);
	MAXIGP0AWQOS			=> open,		-- out std_logic_vector(3 downto 0);
	MAXIGP0AWSIZE			=> open,		-- out std_logic_vector(1 downto 0);
	MAXIGP0AWVALID			=> open,		-- out std_ulogic;
	MAXIGP0BREADY			=> open,		-- out std_ulogic;
	MAXIGP0RREADY			=> open,		-- out std_ulogic;
	MAXIGP0WDATA			=> open,		-- out std_logic_vector(31 downto 0);
	MAXIGP0WID			=> open,		-- out std_logic_vector(11 downto 0);
	MAXIGP0WLAST			=> open,		-- out std_ulogic;
	MAXIGP0WSTRB			=> open,		-- out std_logic_vector(3 downto 0);
	MAXIGP0WVALID			=> open,		-- out std_ulogic;
	MAXIGP1ARADDR			=> open,		-- out std_logic_vector(31 downto 0);
	MAXIGP1ARBURST			=> open,		-- out std_logic_vector(1 downto 0);
	MAXIGP1ARCACHE			=> open,		-- out std_logic_vector(3 downto 0);
	MAXIGP1ARESETN			=> open,		-- out std_ulogic;
	MAXIGP1ARID			=> open,		-- out std_logic_vector(11 downto 0);
	MAXIGP1ARLEN			=> open,		-- out std_logic_vector(3 downto 0);
	MAXIGP1ARLOCK			=> open,		-- out std_logic_vector(1 downto 0);
	MAXIGP1ARPROT			=> open,		-- out std_logic_vector(2 downto 0);
	MAXIGP1ARQOS			=> open,		-- out std_logic_vector(3 downto 0);
	MAXIGP1ARSIZE			=> open,		-- out std_logic_vector(1 downto 0);
	MAXIGP1ARVALID			=> open,		-- out std_ulogic;
	MAXIGP1AWADDR			=> open,		-- out std_logic_vector(31 downto 0);
	MAXIGP1AWBURST			=> open,		-- out std_logic_vector(1 downto 0);
	MAXIGP1AWCACHE			=> open,		-- out std_logic_vector(3 downto 0);
	MAXIGP1AWID			=> open,		-- out std_logic_vector(11 downto 0);
	MAXIGP1AWLEN			=> open,		-- out std_logic_vector(3 downto 0);
	MAXIGP1AWLOCK			=> open,		-- out std_logic_vector(1 downto 0);
	MAXIGP1AWPROT			=> open,		-- out std_logic_vector(2 downto 0);
	MAXIGP1AWQOS			=> open,		-- out std_logic_vector(3 downto 0);
	MAXIGP1AWSIZE			=> open,		-- out std_logic_vector(1 downto 0);
	MAXIGP1AWVALID			=> open,		-- out std_ulogic;
	MAXIGP1BREADY			=> open,		-- out std_ulogic;
	MAXIGP1RREADY			=> open,		-- out std_ulogic;
	MAXIGP1WDATA			=> open,		-- out std_logic_vector(31 downto 0);
	MAXIGP1WID			=> open,		-- out std_logic_vector(11 downto 0);
	MAXIGP1WLAST			=> open,		-- out std_ulogic;
	MAXIGP1WSTRB			=> open,		-- out std_logic_vector(3 downto 0);
	MAXIGP1WVALID			=> open,		-- out std_ulogic;
	SAXIACPARESETN			=> open,		-- out std_ulogic;
	SAXIACPARREADY			=> open,		-- out std_ulogic;
	SAXIACPAWREADY			=> open,		-- out std_ulogic;
	SAXIACPBID			=> open,		-- out std_logic_vector(2 downto 0);
	SAXIACPBRESP			=> open,		-- out std_logic_vector(1 downto 0);
	SAXIACPBVALID			=> open,		-- out std_ulogic;
	SAXIACPRDATA			=> open,		-- out std_logic_vector(63 downto 0);
	SAXIACPRID			=> open,		-- out std_logic_vector(2 downto 0);
	SAXIACPRLAST			=> open,		-- out std_ulogic;
	SAXIACPRRESP			=> open,		-- out std_logic_vector(1 downto 0);
	SAXIACPRVALID			=> open,		-- out std_ulogic;
	SAXIACPWREADY			=> open,		-- out std_ulogic;
	SAXIGP0ARESETN			=> open,		-- out std_ulogic;
	SAXIGP0ARREADY			=> open,		-- out std_ulogic;
	SAXIGP0AWREADY			=> open,		-- out std_ulogic;
	SAXIGP0BID			=> open,		-- out std_logic_vector(5 downto 0);
	SAXIGP0BRESP			=> open,		-- out std_logic_vector(1 downto 0);
	SAXIGP0BVALID			=> open,		-- out std_ulogic;
	SAXIGP0RDATA			=> open,		-- out std_logic_vector(31 downto 0);
	SAXIGP0RID			=> open,		-- out std_logic_vector(5 downto 0);
	SAXIGP0RLAST			=> open,		-- out std_ulogic;
	SAXIGP0RRESP			=> open,		-- out std_logic_vector(1 downto 0);
	SAXIGP0RVALID			=> open,		-- out std_ulogic;
	SAXIGP0WREADY			=> open,		-- out std_ulogic;
	SAXIGP1ARESETN			=> open,		-- out std_ulogic;
	SAXIGP1ARREADY			=> open,		-- out std_ulogic;
	SAXIGP1AWREADY			=> open,		-- out std_ulogic;
	SAXIGP1BID			=> open,		-- out std_logic_vector(5 downto 0);
	SAXIGP1BRESP			=> open,		-- out std_logic_vector(1 downto 0);
	SAXIGP1BVALID			=> open,		-- out std_ulogic;
	SAXIGP1RDATA			=> open,		-- out std_logic_vector(31 downto 0);
	SAXIGP1RID			=> open,		-- out std_logic_vector(5 downto 0);
	SAXIGP1RLAST			=> open,		-- out std_ulogic;
	SAXIGP1RRESP			=> open,		-- out std_logic_vector(1 downto 0);
	SAXIGP1RVALID			=> open,		-- out std_ulogic;
	SAXIGP1WREADY			=> open,		-- out std_ulogic;
	SAXIHP0ARESETN			=> open,		-- out std_ulogic;
	SAXIHP0ARREADY			=> open,		-- out std_ulogic;
	SAXIHP0AWREADY			=> open,		-- out std_ulogic;
	SAXIHP0BID			=> open,		-- out std_logic_vector(5 downto 0);
	SAXIHP0BRESP			=> open,		-- out std_logic_vector(1 downto 0);
	SAXIHP0BVALID			=> open,		-- out std_ulogic;
	SAXIHP0RACOUNT			=> open,		-- out std_logic_vector(2 downto 0);
	SAXIHP0RCOUNT			=> open,		-- out std_logic_vector(7 downto 0);
	SAXIHP0RDATA			=> open,		-- out std_logic_vector(63 downto 0);
	SAXIHP0RID			=> open,		-- out std_logic_vector(5 downto 0);
	SAXIHP0RLAST			=> open,		-- out std_ulogic;
	SAXIHP0RRESP			=> open,		-- out std_logic_vector(1 downto 0);
	SAXIHP0RVALID			=> open,		-- out std_ulogic;
	SAXIHP0WACOUNT			=> open,		-- out std_logic_vector(5 downto 0);
	SAXIHP0WCOUNT			=> open,		-- out std_logic_vector(7 downto 0);
	SAXIHP0WREADY			=> open,		-- out std_ulogic;
	SAXIHP1ARESETN			=> open,		-- out std_ulogic;
	SAXIHP1ARREADY			=> open,		-- out std_ulogic;
	SAXIHP1AWREADY			=> open,		-- out std_ulogic;
	SAXIHP1BID			=> open,		-- out std_logic_vector(5 downto 0);
	SAXIHP1BRESP			=> open,		-- out std_logic_vector(1 downto 0);
	SAXIHP1BVALID			=> open,		-- out std_ulogic;
	SAXIHP1RACOUNT			=> open,		-- out std_logic_vector(2 downto 0);
	SAXIHP1RCOUNT			=> open,		-- out std_logic_vector(7 downto 0);
	SAXIHP1RDATA			=> open,		-- out std_logic_vector(63 downto 0);
	SAXIHP1RID			=> open,		-- out std_logic_vector(5 downto 0);
	SAXIHP1RLAST			=> open,		-- out std_ulogic;
	SAXIHP1RRESP			=> open,		-- out std_logic_vector(1 downto 0);
	SAXIHP1RVALID			=> open,		-- out std_ulogic;
	SAXIHP1WACOUNT			=> open,		-- out std_logic_vector(5 downto 0);
	SAXIHP1WCOUNT			=> open,		-- out std_logic_vector(7 downto 0);
	SAXIHP1WREADY			=> open,		-- out std_ulogic;
	SAXIHP2ARESETN			=> open,		-- out std_ulogic;
	SAXIHP2ARREADY			=> open,		-- out std_ulogic;
	SAXIHP2AWREADY			=> open,		-- out std_ulogic;
	SAXIHP2BID			=> open,		-- out std_logic_vector(5 downto 0);
	SAXIHP2BRESP			=> open,		-- out std_logic_vector(1 downto 0);
	SAXIHP2BVALID			=> open,		-- out std_ulogic;
	SAXIHP2RACOUNT			=> open,		-- out std_logic_vector(2 downto 0);
	SAXIHP2RCOUNT			=> open,		-- out std_logic_vector(7 downto 0);
	SAXIHP2RDATA			=> open,		-- out std_logic_vector(63 downto 0);
	SAXIHP2RID			=> open,		-- out std_logic_vector(5 downto 0);
	SAXIHP2RLAST			=> open,		-- out std_ulogic;
	SAXIHP2RRESP			=> open,		-- out std_logic_vector(1 downto 0);
	SAXIHP2RVALID			=> open,		-- out std_ulogic;
	SAXIHP2WACOUNT			=> open,		-- out std_logic_vector(5 downto 0);
	SAXIHP2WCOUNT			=> open,		-- out std_logic_vector(7 downto 0);
	SAXIHP2WREADY			=> open,		-- out std_ulogic;
	SAXIHP3ARESETN			=> open,		-- out std_ulogic;
	SAXIHP3ARREADY			=> open,		-- out std_ulogic;
	SAXIHP3AWREADY			=> open,		-- out std_ulogic;
	SAXIHP3BID			=> open,		-- out std_logic_vector(5 downto 0);
	SAXIHP3BRESP			=> open,		-- out std_logic_vector(1 downto 0);
	SAXIHP3BVALID			=> open,		-- out std_ulogic;
	SAXIHP3RACOUNT			=> open,		-- out std_logic_vector(2 downto 0);
	SAXIHP3RCOUNT			=> open,		-- out std_logic_vector(7 downto 0);
	SAXIHP3RDATA			=> open,		-- out std_logic_vector(63 downto 0);
	SAXIHP3RID			=> open,		-- out std_logic_vector(5 downto 0);
	SAXIHP3RLAST			=> open,		-- out std_ulogic;
	SAXIHP3RRESP			=> open,		-- out std_logic_vector(1 downto 0);
	SAXIHP3RVALID			=> open,		-- out std_ulogic;
	SAXIHP3WACOUNT			=> open,		-- out std_logic_vector(5 downto 0);
	SAXIHP3WCOUNT			=> open,		-- out std_logic_vector(7 downto 0);
	SAXIHP3WREADY			=> open,		-- out std_ulogic;
	DDRA				=> open,		-- inout std_logic_vector(14 downto 0);
	DDRBA				=> open,		-- inout std_logic_vector(2 downto 0);
	DDRCASB				=> open,		-- inout std_ulogic;
	DDRCKE				=> open,		-- inout std_ulogic;
	DDRCKN				=> open,		-- inout std_ulogic;
	DDRCKP				=> open,		-- inout std_ulogic;
	DDRCSB				=> open,		-- inout std_ulogic;
	DDRDM				=> open,		-- inout std_logic_vector(3 downto 0);
	DDRDQ				=> open,		-- inout std_logic_vector(31 downto 0);
	DDRDQSN				=> open,		-- inout std_logic_vector(3 downto 0);
	DDRDQSP				=> open,		-- inout std_logic_vector(3 downto 0);
	DDRDRSTB			=> open,		-- inout std_ulogic;
	DDRODT				=> open,		-- inout std_ulogic;
	DDRRASB				=> open,		-- inout std_ulogic;
	DDRVRN				=> open,		-- inout std_ulogic;
	DDRVRP				=> open,		-- inout std_ulogic;
	DDRWEB				=> open,		-- inout std_ulogic;
	MIO				=> open,		-- inout std_logic_vector(53 downto 0);
	PSCLK				=> open,		-- inout std_ulogic;
	PSPORB				=> open,		-- inout std_ulogic;
	PSSRSTB				=> open,		-- inout std_ulogic;
	DDRARB				=> (others => '0'),	-- in std_logic_vector(3 downto 0);
	DMA0ACLK			=> '0', 		-- in std_ulogic;
	DMA0DAREADY			=> '0', 		-- in std_ulogic;
	DMA0DRLAST			=> '0', 		-- in std_ulogic;
	DMA0DRTYPE			=> (others => '0'),	-- in std_logic_vector(1 downto 0);
	DMA0DRVALID			=> '0', 		-- in std_ulogic;
	DMA1ACLK			=> '0', 		-- in std_ulogic;
	DMA1DAREADY			=> '0', 		-- in std_ulogic;
	DMA1DRLAST			=> '0', 		-- in std_ulogic;
	DMA1DRTYPE			=> (others => '0'),	-- in std_logic_vector(1 downto 0);
	DMA1DRVALID			=> '0', 		-- in std_ulogic;
	DMA2ACLK			=> '0', 		-- in std_ulogic;
	DMA2DAREADY			=> '0', 		-- in std_ulogic;
	DMA2DRLAST			=> '0', 		-- in std_ulogic;
	DMA2DRTYPE			=> (others => '0'),	-- in std_logic_vector(1 downto 0);
	DMA2DRVALID			=> '0', 		-- in std_ulogic;
	DMA3ACLK			=> '0', 		-- in std_ulogic;
	DMA3DAREADY			=> '0', 		-- in std_ulogic;
	DMA3DRLAST			=> '0', 		-- in std_ulogic;
	DMA3DRTYPE			=> (others => '0'),	-- in std_logic_vector(1 downto 0);
	DMA3DRVALID			=> '0', 		-- in std_ulogic;
	EMIOCAN0PHYRX			=> '0', 		-- in std_ulogic;
	EMIOCAN1PHYRX			=> '0', 		-- in std_ulogic;
	EMIOENET0EXTINTIN		=> '0', 		-- in std_ulogic;
	EMIOENET0GMIICOL		=> '0', 		-- in std_ulogic;
	EMIOENET0GMIICRS		=> '0', 		-- in std_ulogic;
	EMIOENET0GMIIRXCLK		=> '0', 		-- in std_ulogic;
	EMIOENET0GMIIRXD		=> (others => '0'),	-- in std_logic_vector(7 downto 0);
	EMIOENET0GMIIRXDV		=> '0', 		-- in std_ulogic;
	EMIOENET0GMIIRXER		=> '0', 		-- in std_ulogic;
	EMIOENET0GMIITXCLK		=> '0', 		-- in std_ulogic;
	EMIOENET0MDIOI			=> '0', 		-- in std_ulogic;
	EMIOENET1EXTINTIN		=> '0', 		-- in std_ulogic;
	EMIOENET1GMIICOL		=> '0', 		-- in std_ulogic;
	EMIOENET1GMIICRS		=> '0', 		-- in std_ulogic;
	EMIOENET1GMIIRXCLK		=> '0', 		-- in std_ulogic;
	EMIOENET1GMIIRXD		=> (others => '0'),	-- in std_logic_vector(7 downto 0);
	EMIOENET1GMIIRXDV		=> '0', 		-- in std_ulogic;
	EMIOENET1GMIIRXER		=> '0', 		-- in std_ulogic;
	EMIOENET1GMIITXCLK		=> '0', 		-- in std_ulogic;
	EMIOENET1MDIOI			=> '0', 		-- in std_ulogic;
	EMIOGPIOI			=> (others => '0'),	-- in std_logic_vector(63 downto 0);
	EMIOI2C0SCLI			=> '0', 		-- in std_ulogic;
	EMIOI2C0SDAI			=> '0', 		-- in std_ulogic;
	EMIOI2C1SCLI			=> '0', 		-- in std_ulogic;
	EMIOI2C1SDAI			=> '0', 		-- in std_ulogic;
	EMIOPJTAGTCK			=> '0', 		-- in std_ulogic;
	EMIOPJTAGTDI			=> '0', 		-- in std_ulogic;
	EMIOPJTAGTMS			=> '0', 		-- in std_ulogic;
	EMIOSDIO0CDN			=> '0', 		-- in std_ulogic;
	EMIOSDIO0CLKFB			=> '0', 		-- in std_ulogic;
	EMIOSDIO0CMDI			=> '0', 		-- in std_ulogic;
	EMIOSDIO0DATAI			=> (others => '0'),	-- in std_logic_vector(3 downto 0);
	EMIOSDIO0WP			=> '0', 		-- in std_ulogic;
	EMIOSDIO1CDN			=> '0', 		-- in std_ulogic;
	EMIOSDIO1CLKFB			=> '0', 		-- in std_ulogic;
	EMIOSDIO1CMDI			=> '0', 		-- in std_ulogic;
	EMIOSDIO1DATAI			=> (others => '0'),	-- in std_logic_vector(3 downto 0);
	EMIOSDIO1WP			=> '0', 		-- in std_ulogic;
	EMIOSPI0MI			=> '0', 		-- in std_ulogic;
	EMIOSPI0SCLKI			=> '0', 		-- in std_ulogic;
	EMIOSPI0SI			=> '0', 		-- in std_ulogic;
	EMIOSPI0SSIN			=> '0', 		-- in std_ulogic;
	EMIOSPI1MI			=> '0', 		-- in std_ulogic;
	EMIOSPI1SCLKI			=> '0', 		-- in std_ulogic;
	EMIOSPI1SI			=> '0', 		-- in std_ulogic;
	EMIOSPI1SSIN			=> '0', 		-- in std_ulogic;
	EMIOSRAMINTIN			=> '0', 		-- in std_ulogic;
	EMIOTRACECLK			=> '0', 		-- in std_ulogic;
	EMIOTTC0CLKI			=> (others => '0'),	-- in std_logic_vector(2 downto 0);
	EMIOTTC1CLKI			=> (others => '0'),	-- in std_logic_vector(2 downto 0);
	EMIOUART0CTSN			=> '0', 		-- in std_ulogic;
	EMIOUART0DCDN			=> '0', 		-- in std_ulogic;
	EMIOUART0DSRN			=> '0', 		-- in std_ulogic;
	EMIOUART0RIN			=> '0', 		-- in std_ulogic;
	EMIOUART0RX			=> '0', 		-- in std_ulogic;
	EMIOUART1CTSN			=> '0', 		-- in std_ulogic;
	EMIOUART1DCDN			=> '0', 		-- in std_ulogic;
	EMIOUART1DSRN			=> '0', 		-- in std_ulogic;
	EMIOUART1RIN			=> '0', 		-- in std_ulogic;
	EMIOUART1RX			=> '0', 		-- in std_ulogic;
	EMIOUSB0VBUSPWRFAULT		=> '0', 		-- in std_ulogic;
	EMIOUSB1VBUSPWRFAULT		=> '0', 		-- in std_ulogic;
	EMIOWDTCLKI			=> '0', 		-- in std_ulogic;
	EVENTEVENTI			=> '0', 		-- in std_ulogic;
	FCLKCLKTRIGN			=> (others => '0'),	-- in std_logic_vector(3 downto 0);
	FPGAIDLEN			=> '0', 		-- in std_ulogic;
	FTMDTRACEINATID			=> (others => '0'),	-- in std_logic_vector(3 downto 0);
	FTMDTRACEINCLOCK		=> '0', 		-- in std_ulogic;
	FTMDTRACEINDATA			=> (others => '0'),	-- in std_logic_vector(31 downto 0);
	FTMDTRACEINVALID		=> '0', 		-- in std_ulogic;
	FTMTF2PDEBUG			=> (others => '0'),	-- in std_logic_vector(31 downto 0);
	FTMTF2PTRIG			=> (others => '0'),	-- in std_logic_vector(3 downto 0);
	FTMTP2FTRIGACK			=> (others => '0'),	-- in std_logic_vector(3 downto 0);
	IRQF2P				=> (others => '0'),	-- in std_logic_vector(19 downto 0);
	MAXIGP0ACLK			=> '0', 		-- in std_ulogic;
	MAXIGP0ARREADY			=> '0', 		-- in std_ulogic;
	MAXIGP0AWREADY			=> '0', 		-- in std_ulogic;
	MAXIGP0BID			=> (others => '0'),	-- in std_logic_vector(11 downto 0);
	MAXIGP0BRESP			=> (others => '0'),	-- in std_logic_vector(1 downto 0);
	MAXIGP0BVALID			=> '0', 		-- in std_ulogic;
	MAXIGP0RDATA			=> (others => '0'),	-- in std_logic_vector(31 downto 0);
	MAXIGP0RID			=> (others => '0'),	-- in std_logic_vector(11 downto 0);
	MAXIGP0RLAST			=> '0', 		-- in std_ulogic;
	MAXIGP0RRESP			=> (others => '0'),	-- in std_logic_vector(1 downto 0);
	MAXIGP0RVALID			=> '0', 		-- in std_ulogic;
	MAXIGP0WREADY			=> '0', 		-- in std_ulogic;
	MAXIGP1ACLK			=> '0', 		-- in std_ulogic;
	MAXIGP1ARREADY			=> '0', 		-- in std_ulogic;
	MAXIGP1AWREADY			=> '0', 		-- in std_ulogic;
	MAXIGP1BID			=> (others => '0'),	-- in std_logic_vector(11 downto 0);
	MAXIGP1BRESP			=> (others => '0'),	-- in std_logic_vector(1 downto 0);
	MAXIGP1BVALID			=> '0', 		-- in std_ulogic;
	MAXIGP1RDATA			=> (others => '0'),	-- in std_logic_vector(31 downto 0);
	MAXIGP1RID			=> (others => '0'),	-- in std_logic_vector(11 downto 0);
	MAXIGP1RLAST			=> '0', 		-- in std_ulogic;
	MAXIGP1RRESP			=> (others => '0'),	-- in std_logic_vector(1 downto 0);
	MAXIGP1RVALID			=> '0', 		-- in std_ulogic;
	MAXIGP1WREADY			=> '0', 		-- in std_ulogic;
	SAXIACPACLK			=> '0', 		-- in std_ulogic;
	SAXIACPARADDR			=> (others => '0'),	-- in std_logic_vector(31 downto 0);
	SAXIACPARBURST			=> (others => '0'),	-- in std_logic_vector(1 downto 0);
	SAXIACPARCACHE			=> (others => '0'),	-- in std_logic_vector(3 downto 0);
	SAXIACPARID			=> (others => '0'),	-- in std_logic_vector(2 downto 0);
	SAXIACPARLEN			=> (others => '0'),	-- in std_logic_vector(3 downto 0);
	SAXIACPARLOCK			=> (others => '0'),	-- in std_logic_vector(1 downto 0);
	SAXIACPARPROT			=> (others => '0'),	-- in std_logic_vector(2 downto 0);
	SAXIACPARQOS			=> (others => '0'),	-- in std_logic_vector(3 downto 0);
	SAXIACPARSIZE			=> (others => '0'),	-- in std_logic_vector(1 downto 0);
	SAXIACPARUSER			=> (others => '0'),	-- in std_logic_vector(4 downto 0);
	SAXIACPARVALID			=> '0', 		-- in std_ulogic;
	SAXIACPAWADDR			=> (others => '0'),	-- in std_logic_vector(31 downto 0);
	SAXIACPAWBURST			=> (others => '0'),	-- in std_logic_vector(1 downto 0);
	SAXIACPAWCACHE			=> (others => '0'),	-- in std_logic_vector(3 downto 0);
	SAXIACPAWID			=> (others => '0'),	-- in std_logic_vector(2 downto 0);
	SAXIACPAWLEN			=> (others => '0'),	-- in std_logic_vector(3 downto 0);
	SAXIACPAWLOCK			=> (others => '0'),	-- in std_logic_vector(1 downto 0);
	SAXIACPAWPROT			=> (others => '0'),	-- in std_logic_vector(2 downto 0);
	SAXIACPAWQOS			=> (others => '0'),	-- in std_logic_vector(3 downto 0);
	SAXIACPAWSIZE			=> (others => '0'),	-- in std_logic_vector(1 downto 0);
	SAXIACPAWUSER			=> (others => '0'),	-- in std_logic_vector(4 downto 0);
	SAXIACPAWVALID			=> '0', 		-- in std_ulogic;
	SAXIACPBREADY			=> '0', 		-- in std_ulogic;
	SAXIACPRREADY			=> '0', 		-- in std_ulogic;
	SAXIACPWDATA			=> (others => '0'),	-- in std_logic_vector(63 downto 0);
	SAXIACPWID			=> (others => '0'),	-- in std_logic_vector(2 downto 0);
	SAXIACPWLAST			=> '0', 		-- in std_ulogic;
	SAXIACPWSTRB			=> (others => '0'),	-- in std_logic_vector(7 downto 0);
	SAXIACPWVALID			=> '0', 		-- in std_ulogic;
	SAXIGP0ACLK			=> '0', 		-- in std_ulogic;
	SAXIGP0ARADDR			=> (others => '0'),	-- in std_logic_vector(31 downto 0);
	SAXIGP0ARBURST			=> (others => '0'),	-- in std_logic_vector(1 downto 0);
	SAXIGP0ARCACHE			=> (others => '0'),	-- in std_logic_vector(3 downto 0);
	SAXIGP0ARID			=> (others => '0'),	-- in std_logic_vector(5 downto 0);
	SAXIGP0ARLEN			=> (others => '0'),	-- in std_logic_vector(3 downto 0);
	SAXIGP0ARLOCK			=> (others => '0'),	-- in std_logic_vector(1 downto 0);
	SAXIGP0ARPROT			=> (others => '0'),	-- in std_logic_vector(2 downto 0);
	SAXIGP0ARQOS			=> (others => '0'),	-- in std_logic_vector(3 downto 0);
	SAXIGP0ARSIZE			=> (others => '0'),	-- in std_logic_vector(1 downto 0);
	SAXIGP0ARVALID			=> '0', 		-- in std_ulogic;
	SAXIGP0AWADDR			=> (others => '0'),	-- in std_logic_vector(31 downto 0);
	SAXIGP0AWBURST			=> (others => '0'),	-- in std_logic_vector(1 downto 0);
	SAXIGP0AWCACHE			=> (others => '0'),	-- in std_logic_vector(3 downto 0);
	SAXIGP0AWID			=> (others => '0'),	-- in std_logic_vector(5 downto 0);
	SAXIGP0AWLEN			=> (others => '0'),	-- in std_logic_vector(3 downto 0);
	SAXIGP0AWLOCK			=> (others => '0'),	-- in std_logic_vector(1 downto 0);
	SAXIGP0AWPROT			=> (others => '0'),	-- in std_logic_vector(2 downto 0);
	SAXIGP0AWQOS			=> (others => '0'),	-- in std_logic_vector(3 downto 0);
	SAXIGP0AWSIZE			=> (others => '0'),	-- in std_logic_vector(1 downto 0);
	SAXIGP0AWVALID			=> '0', 		-- in std_ulogic;
	SAXIGP0BREADY			=> '0', 		-- in std_ulogic;
	SAXIGP0RREADY			=> '0', 		-- in std_ulogic;
	SAXIGP0WDATA			=> (others => '0'),	-- in std_logic_vector(31 downto 0);
	SAXIGP0WID			=> (others => '0'),	-- in std_logic_vector(5 downto 0);
	SAXIGP0WLAST			=> '0', 		-- in std_ulogic;
	SAXIGP0WSTRB			=> (others => '0'),	-- in std_logic_vector(3 downto 0);
	SAXIGP0WVALID			=> '0', 		-- in std_ulogic;
	SAXIGP1ACLK			=> '0', 		-- in std_ulogic;
	SAXIGP1ARADDR			=> (others => '0'),	-- in std_logic_vector(31 downto 0);
	SAXIGP1ARBURST			=> (others => '0'),	-- in std_logic_vector(1 downto 0);
	SAXIGP1ARCACHE			=> (others => '0'),	-- in std_logic_vector(3 downto 0);
	SAXIGP1ARID			=> (others => '0'),	-- in std_logic_vector(5 downto 0);
	SAXIGP1ARLEN			=> (others => '0'),	-- in std_logic_vector(3 downto 0);
	SAXIGP1ARLOCK			=> (others => '0'),	-- in std_logic_vector(1 downto 0);
	SAXIGP1ARPROT			=> (others => '0'),	-- in std_logic_vector(2 downto 0);
	SAXIGP1ARQOS			=> (others => '0'),	-- in std_logic_vector(3 downto 0);
	SAXIGP1ARSIZE			=> (others => '0'),	-- in std_logic_vector(1 downto 0);
	SAXIGP1ARVALID			=> '0', 		-- in std_ulogic;
	SAXIGP1AWADDR			=> (others => '0'),	-- in std_logic_vector(31 downto 0);
	SAXIGP1AWBURST			=> (others => '0'),	-- in std_logic_vector(1 downto 0);
	SAXIGP1AWCACHE			=> (others => '0'),	-- in std_logic_vector(3 downto 0);
	SAXIGP1AWID			=> (others => '0'),	-- in std_logic_vector(5 downto 0);
	SAXIGP1AWLEN			=> (others => '0'),	-- in std_logic_vector(3 downto 0);
	SAXIGP1AWLOCK			=> (others => '0'),	-- in std_logic_vector(1 downto 0);
	SAXIGP1AWPROT			=> (others => '0'),	-- in std_logic_vector(2 downto 0);
	SAXIGP1AWQOS			=> (others => '0'),	-- in std_logic_vector(3 downto 0);
	SAXIGP1AWSIZE			=> (others => '0'),	-- in std_logic_vector(1 downto 0);
	SAXIGP1AWVALID			=> '0', 		-- in std_ulogic;
	SAXIGP1BREADY			=> '0', 		-- in std_ulogic;
	SAXIGP1RREADY			=> '0', 		-- in std_ulogic;
	SAXIGP1WDATA			=> (others => '0'),	-- in std_logic_vector(31 downto 0);
	SAXIGP1WID			=> (others => '0'),	-- in std_logic_vector(5 downto 0);
	SAXIGP1WLAST			=> '0', 		-- in std_ulogic;
	SAXIGP1WSTRB			=> (others => '0'),	-- in std_logic_vector(3 downto 0);
	SAXIGP1WVALID			=> '0', 		-- in std_ulogic;
	SAXIHP0ACLK			=> '0', 		-- in std_ulogic;
	SAXIHP0ARADDR			=> (others => '0'),	-- in std_logic_vector(31 downto 0);
	SAXIHP0ARBURST			=> (others => '0'),	-- in std_logic_vector(1 downto 0);
	SAXIHP0ARCACHE			=> (others => '0'),	-- in std_logic_vector(3 downto 0);
	SAXIHP0ARID			=> (others => '0'),	-- in std_logic_vector(5 downto 0);
	SAXIHP0ARLEN			=> (others => '0'),	-- in std_logic_vector(3 downto 0);
	SAXIHP0ARLOCK			=> (others => '0'),	-- in std_logic_vector(1 downto 0);
	SAXIHP0ARPROT			=> (others => '0'),	-- in std_logic_vector(2 downto 0);
	SAXIHP0ARQOS			=> (others => '0'),	-- in std_logic_vector(3 downto 0);
	SAXIHP0ARSIZE			=> (others => '0'),	-- in std_logic_vector(1 downto 0);
	SAXIHP0ARVALID			=> '0', 		-- in std_ulogic;
	SAXIHP0AWADDR			=> (others => '0'),	-- in std_logic_vector(31 downto 0);
	SAXIHP0AWBURST			=> (others => '0'),	-- in std_logic_vector(1 downto 0);
	SAXIHP0AWCACHE			=> (others => '0'),	-- in std_logic_vector(3 downto 0);
	SAXIHP0AWID			=> (others => '0'),	-- in std_logic_vector(5 downto 0);
	SAXIHP0AWLEN			=> (others => '0'),	-- in std_logic_vector(3 downto 0);
	SAXIHP0AWLOCK			=> (others => '0'),	-- in std_logic_vector(1 downto 0);
	SAXIHP0AWPROT			=> (others => '0'),	-- in std_logic_vector(2 downto 0);
	SAXIHP0AWQOS			=> (others => '0'),	-- in std_logic_vector(3 downto 0);
	SAXIHP0AWSIZE			=> (others => '0'),	-- in std_logic_vector(1 downto 0);
	SAXIHP0AWVALID			=> '0', 		-- in std_ulogic;
	SAXIHP0BREADY			=> '0', 		-- in std_ulogic;
	SAXIHP0RDISSUECAP1EN		=> '0', 		-- in std_ulogic;
	SAXIHP0RREADY			=> '0', 		-- in std_ulogic;
	SAXIHP0WDATA			=> (others => '0'),	-- in std_logic_vector(63 downto 0);
	SAXIHP0WID			=> (others => '0'),	-- in std_logic_vector(5 downto 0);
	SAXIHP0WLAST			=> '0', 		-- in std_ulogic;
	SAXIHP0WRISSUECAP1EN		=> '0', 		-- in std_ulogic;
	SAXIHP0WSTRB			=> (others => '0'),	-- in std_logic_vector(7 downto 0);
	SAXIHP0WVALID			=> '0', 		-- in std_ulogic;
	SAXIHP1ACLK			=> '0', 		-- in std_ulogic;
	SAXIHP1ARADDR			=> (others => '0'),	-- in std_logic_vector(31 downto 0);
	SAXIHP1ARBURST			=> (others => '0'),	-- in std_logic_vector(1 downto 0);
	SAXIHP1ARCACHE			=> (others => '0'),	-- in std_logic_vector(3 downto 0);
	SAXIHP1ARID			=> (others => '0'),	-- in std_logic_vector(5 downto 0);
	SAXIHP1ARLEN			=> (others => '0'),	-- in std_logic_vector(3 downto 0);
	SAXIHP1ARLOCK			=> (others => '0'),	-- in std_logic_vector(1 downto 0);
	SAXIHP1ARPROT			=> (others => '0'),	-- in std_logic_vector(2 downto 0);
	SAXIHP1ARQOS			=> (others => '0'),	-- in std_logic_vector(3 downto 0);
	SAXIHP1ARSIZE			=> (others => '0'),	-- in std_logic_vector(1 downto 0);
	SAXIHP1ARVALID			=> '0', 		-- in std_ulogic;
	SAXIHP1AWADDR			=> (others => '0'),	-- in std_logic_vector(31 downto 0);
	SAXIHP1AWBURST			=> (others => '0'),	-- in std_logic_vector(1 downto 0);
	SAXIHP1AWCACHE			=> (others => '0'),	-- in std_logic_vector(3 downto 0);
	SAXIHP1AWID			=> (others => '0'),	-- in std_logic_vector(5 downto 0);
	SAXIHP1AWLEN			=> (others => '0'),	-- in std_logic_vector(3 downto 0);
	SAXIHP1AWLOCK			=> (others => '0'),	-- in std_logic_vector(1 downto 0);
	SAXIHP1AWPROT			=> (others => '0'),	-- in std_logic_vector(2 downto 0);
	SAXIHP1AWQOS			=> (others => '0'),	-- in std_logic_vector(3 downto 0);
	SAXIHP1AWSIZE			=> (others => '0'),	-- in std_logic_vector(1 downto 0);
	SAXIHP1AWVALID			=> '0', 		-- in std_ulogic;
	SAXIHP1BREADY			=> '0', 		-- in std_ulogic;
	SAXIHP1RDISSUECAP1EN		=> '0', 		-- in std_ulogic;
	SAXIHP1RREADY			=> '0', 		-- in std_ulogic;
	SAXIHP1WDATA			=> (others => '0'),	-- in std_logic_vector(63 downto 0);
	SAXIHP1WID			=> (others => '0'),	-- in std_logic_vector(5 downto 0);
	SAXIHP1WLAST			=> '0', 		-- in std_ulogic;
	SAXIHP1WRISSUECAP1EN		=> '0', 		-- in std_ulogic;
	SAXIHP1WSTRB			=> (others => '0'),	-- in std_logic_vector(7 downto 0);
	SAXIHP1WVALID			=> '0', 		-- in std_ulogic;
	SAXIHP2ACLK			=> '0', 		-- in std_ulogic;
	SAXIHP2ARADDR			=> (others => '0'),	-- in std_logic_vector(31 downto 0);
	SAXIHP2ARBURST			=> (others => '0'),	-- in std_logic_vector(1 downto 0);
	SAXIHP2ARCACHE			=> (others => '0'),	-- in std_logic_vector(3 downto 0);
	SAXIHP2ARID			=> (others => '0'),	-- in std_logic_vector(5 downto 0);
	SAXIHP2ARLEN			=> (others => '0'),	-- in std_logic_vector(3 downto 0);
	SAXIHP2ARLOCK			=> (others => '0'),	-- in std_logic_vector(1 downto 0);
	SAXIHP2ARPROT			=> (others => '0'),	-- in std_logic_vector(2 downto 0);
	SAXIHP2ARQOS			=> (others => '0'),	-- in std_logic_vector(3 downto 0);
	SAXIHP2ARSIZE			=> (others => '0'),	-- in std_logic_vector(1 downto 0);
	SAXIHP2ARVALID			=> '0', 		-- in std_ulogic;
	SAXIHP2AWADDR			=> (others => '0'),	-- in std_logic_vector(31 downto 0);
	SAXIHP2AWBURST			=> (others => '0'),	-- in std_logic_vector(1 downto 0);
	SAXIHP2AWCACHE			=> (others => '0'),	-- in std_logic_vector(3 downto 0);
	SAXIHP2AWID			=> (others => '0'),	-- in std_logic_vector(5 downto 0);
	SAXIHP2AWLEN			=> (others => '0'),	-- in std_logic_vector(3 downto 0);
	SAXIHP2AWLOCK			=> (others => '0'),	-- in std_logic_vector(1 downto 0);
	SAXIHP2AWPROT			=> (others => '0'),	-- in std_logic_vector(2 downto 0);
	SAXIHP2AWQOS			=> (others => '0'),	-- in std_logic_vector(3 downto 0);
	SAXIHP2AWSIZE			=> (others => '0'),	-- in std_logic_vector(1 downto 0);
	SAXIHP2AWVALID			=> '0', 		-- in std_ulogic;
	SAXIHP2BREADY			=> '0', 		-- in std_ulogic;
	SAXIHP2RDISSUECAP1EN		=> '0', 		-- in std_ulogic;
	SAXIHP2RREADY			=> '0', 		-- in std_ulogic;
	SAXIHP2WDATA			=> (others => '0'),	-- in std_logic_vector(63 downto 0);
	SAXIHP2WID			=> (others => '0'),	-- in std_logic_vector(5 downto 0);
	SAXIHP2WLAST			=> '0', 		-- in std_ulogic;
	SAXIHP2WRISSUECAP1EN		=> '0', 		-- in std_ulogic;
	SAXIHP2WSTRB			=> (others => '0'),	-- in std_logic_vector(7 downto 0);
	SAXIHP2WVALID			=> '0', 		-- in std_ulogic;
	SAXIHP3ACLK			=> '0', 		-- in std_ulogic;
	SAXIHP3ARADDR			=> (others => '0'),	-- in std_logic_vector(31 downto 0);
	SAXIHP3ARBURST			=> (others => '0'),	-- in std_logic_vector(1 downto 0);
	SAXIHP3ARCACHE			=> (others => '0'),	-- in std_logic_vector(3 downto 0);
	SAXIHP3ARID			=> (others => '0'),	-- in std_logic_vector(5 downto 0);
	SAXIHP3ARLEN			=> (others => '0'),	-- in std_logic_vector(3 downto 0);
	SAXIHP3ARLOCK			=> (others => '0'),	-- in std_logic_vector(1 downto 0);
	SAXIHP3ARPROT			=> (others => '0'),	-- in std_logic_vector(2 downto 0);
	SAXIHP3ARQOS			=> (others => '0'),	-- in std_logic_vector(3 downto 0);
	SAXIHP3ARSIZE			=> (others => '0'),	-- in std_logic_vector(1 downto 0);
	SAXIHP3ARVALID			=> '0', 		-- in std_ulogic;
	SAXIHP3AWADDR			=> (others => '0'),	-- in std_logic_vector(31 downto 0);
	SAXIHP3AWBURST			=> (others => '0'),	-- in std_logic_vector(1 downto 0);
	SAXIHP3AWCACHE			=> (others => '0'),	-- in std_logic_vector(3 downto 0);
	SAXIHP3AWID			=> (others => '0'),	-- in std_logic_vector(5 downto 0);
	SAXIHP3AWLEN			=> (others => '0'),	-- in std_logic_vector(3 downto 0);
	SAXIHP3AWLOCK			=> (others => '0'),	-- in std_logic_vector(1 downto 0);
	SAXIHP3AWPROT			=> (others => '0'),	-- in std_logic_vector(2 downto 0);
	SAXIHP3AWQOS			=> (others => '0'),	-- in std_logic_vector(3 downto 0);
	SAXIHP3AWSIZE			=> (others => '0'),	-- in std_logic_vector(1 downto 0);
	SAXIHP3AWVALID			=> '0', 		-- in std_ulogic;
	SAXIHP3BREADY			=> '0', 		-- in std_ulogic;
	SAXIHP3RDISSUECAP1EN		=> '0', 		-- in std_ulogic;
	SAXIHP3RREADY			=> '0', 		-- in std_ulogic;
	SAXIHP3WDATA			=> (others => '0'),	-- in std_logic_vector(63 downto 0);
	SAXIHP3WID			=> (others => '0'),	-- in std_logic_vector(5 downto 0);
	SAXIHP3WLAST			=> '0', 		-- in std_ulogic;
	SAXIHP3WRISSUECAP1EN		=> '0', 		-- in std_ulogic;
	SAXIHP3WSTRB			=> (others => '0'),	-- in std_logic_vector(7 downto 0);
	SAXIHP3WVALID			=> '0'			-- in std_ulogic
    );
	
  process(sysclk)
  begin
    if rising_edge(sysclk) then
      counter <= counter + 1;
    end if;
  end process;

  led <= std_logic_vector(resize(shift_right(counter, 4 * to_integer(unsigned(sw))), 4));
end behaviour;
