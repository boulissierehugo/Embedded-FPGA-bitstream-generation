LIBRARY ieee;
USE ieee.std_logic_1164.ALL;

ENTITY s_box IS
PORT(
    s_in    :	IN  STD_LOGIC_VECTOR(7 DOWNTO 0);
    s_out   :	OUT STD_LOGIC_VECTOR(7 DOWNTO 0)
    );
END s_box;

ARCHITECTURE beh OF s_box IS
    
BEGIN

process (s_in)
begin 
case s_in is 
	-- first row
	WHEN "00000000" => s_out<= "01100011";
	WHEN "00000001" => s_out<= "01111100";
	WHEN "00000010" => s_out<= "01110111";
	WHEN "00000011" => s_out<= "01111011";
	WHEN "00000100" => s_out<= "11110010";
	WHEN "00000101" => s_out<= "01101011";
	WHEN "00000110" => s_out<= "01101111";
	WHEN "00000111" => s_out<= "11000101";
	WHEN "00001000" => s_out<= "00110000";
	WHEN "00001001" => s_out<= "00000001";
	WHEN "00001010" => s_out<= "01100111";
	WHEN "00001011" => s_out<= "00101011";
	WHEN "00001100" => s_out<= "11111110";
	WHEN "00001101" => s_out<= "11010111";
	WHEN "00001110" => s_out<= "10101011";
	WHEN "00001111" => s_out<= "01110110";
	--second row
	WHEN "00010000" => s_out<= "11001010";
	WHEN "00010001" => s_out<= "10000010";
	WHEN "00010010" => s_out<= "11001001";
	WHEN "00010011" => s_out<= "01111101";
	WHEN "00010100" => s_out<= "11111010";
	WHEN "00010101" => s_out<= "01011001";
	WHEN "00010110" => s_out<= "01000111";
	WHEN "00010111" => s_out<= "11110000";
	WHEN "00011000" => s_out<= "10101101";
	WHEN "00011001" => s_out<= "11010100";
	WHEN "00011010" => s_out<= "10100010";
	WHEN "00011011" => s_out<= "10101111";
	WHEN "00011100" => s_out<= "10011100";
	WHEN "00011101" => s_out<= "10100100";
	WHEN "00011110" => s_out<= "01110010";
	WHEN "00011111" => s_out<= "11000000";
	--third row
	WHEN "00100000" => s_out<= "10110111";
	WHEN "00100001" => s_out<= "11111101";
	WHEN "00100010" => s_out<= "10010011";
	WHEN "00100011" => s_out<= "00100110";
	WHEN "00100100" => s_out<= "00110110";
	WHEN "00100101" => s_out<= "00111111";
	WHEN "00100110" => s_out<= "11110111";
	WHEN "00100111" => s_out<= "11001100";
	WHEN "00101000" => s_out<= "00110100";
	WHEN "00101001" => s_out<= "10100101";
	WHEN "00101010" => s_out<= "11100101";
	WHEN "00101011" => s_out<= "11110001";
	WHEN "00101100" => s_out<= "01110001";
	WHEN "00101101" => s_out<= "11011000";
	WHEN "00101110" => s_out<= "00110001";
	WHEN "00101111" => s_out<= "00010101";
	 --forth row
	WHEN "00110000" => s_out<= "00000100";
	WHEN "00110001" => s_out<= "11000111";
	WHEN "00110010" => s_out<= "00100011";
	WHEN "00110011" => s_out<= "11000011";
	WHEN "00110100" => s_out<= "00011000";
	WHEN "00110101" => s_out<= "10010110";
	WHEN "00110110" => s_out<= "00000101";
	WHEN "00110111" => s_out<= "10011010";
	WHEN "00111000" => s_out<= "00000111";
	WHEN "00111001" => s_out<= "00010010";
	WHEN "00111010" => s_out<= "10000000";
	WHEN "00111011" => s_out<= "11100010";
	WHEN "00111100" => s_out<= "11101011";
	WHEN "00111101" => s_out<= "00100111";
	WHEN "00111110" => s_out<= "10110010";
	WHEN "00111111" => s_out<= "01110101";
	--fifth row
	WHEN "01000000" => s_out<= "00001001";
	WHEN "01000001" => s_out<= "10000011";
	WHEN "01000010" => s_out<= "00101100";
	WHEN "01000011" => s_out<= "00011010";
	WHEN "01000100" => s_out<= "00011011";
	WHEN "01000101" => s_out<= "01101110";
	WHEN "01000110" => s_out<= "01011010";
	WHEN "01000111" => s_out<= "10100000";
	WHEN "01001000" => s_out<= "01010010";
	WHEN "01001001" => s_out<= "00111011";
	WHEN "01001010" => s_out<= "11010110";
	WHEN "01001011" => s_out<= "10110011";
	WHEN "01001100" => s_out<= "00101001";
	WHEN "01001101" => s_out<= "11100011";
	WHEN "01001110" => s_out<= "00101111";
	WHEN "01001111" => s_out<= "10000100";
	--sixth row
	WHEN "01010000" => s_out<= "01010011";
	WHEN "01010001" => s_out<= "11010001";
	WHEN "01010010" => s_out<= "00000000";
	WHEN "01010011" => s_out<= "11101101";
	WHEN "01010100" => s_out<= "00100000";
	WHEN "01010101" => s_out<= "11111100";
	WHEN "01010110" => s_out<= "10110001";
	WHEN "01010111" => s_out<= "01011011";
	WHEN "01011000" => s_out<= "01101010";
	WHEN "01011001" => s_out<= "11001011";
	WHEN "01011010" => s_out<= "10111110";
	WHEN "01011011" => s_out<= "00111001";
	WHEN "01011100" => s_out<= "01001010";
	WHEN "01011101" => s_out<= "01001100";
	WHEN "01011110" => s_out<= "01011000";
	WHEN "01011111" => s_out<= "11001111";
	--seventh row	    
	WHEN "01100000" => s_out<= "11010000";
	WHEN "01100001" => s_out<= "11101111";
	WHEN "01100010" => s_out<= "10101010";
	WHEN "01100011" => s_out<= "11111011";
	WHEN "01100100" => s_out<= "01000011";
	WHEN "01100101" => s_out<= "01001101";
	WHEN "01100110" => s_out<= "00110011";
	WHEN "01100111" => s_out<= "10000101";
	WHEN "01101000" => s_out<= "01000101";
	WHEN "01101001" => s_out<= "11111001";
	WHEN "01101010" => s_out<= "00000010";
	WHEN "01101011" => s_out<= "01111111";
	WHEN "01101100" => s_out<= "01010000";
	WHEN "01101101" => s_out<= "00111100";
	WHEN "01101110" => s_out<= "10011111";
	WHEN "01101111" => s_out<= "10101000";
	--eighth row	    
	WHEN "01110000" => s_out<= "01010001";
	WHEN "01110001" => s_out<= "10100011";
	WHEN "01110010" => s_out<= "01000000";
	WHEN "01110011" => s_out<= "10001111";
	WHEN "01110100" => s_out<= "10010010";
	WHEN "01110101" => s_out<= "10011101";
	WHEN "01110110" => s_out<= "00111000";
	WHEN "01110111" => s_out<= "11110101";
	WHEN "01111000" => s_out<= "10111100";
	WHEN "01111001" => s_out<= "10110110";
	WHEN "01111010" => s_out<= "11011010";
	WHEN "01111011" => s_out<= "00100001";
	WHEN "01111100" => s_out<= "00010000";
	WHEN "01111101" => s_out<= "11111111";
	WHEN "01111110" => s_out<= "11110011";
	WHEN "01111111" => s_out<= "11010010";
	--ninth row	  
	WHEN "10000000" => s_out<= "11001101";
	WHEN "10000001" => s_out<= "00001100";
	WHEN "10000010" => s_out<= "00010011";
	WHEN "10000011" => s_out<= "11101100";
	WHEN "10000100" => s_out<= "01011111";
	WHEN "10000101" => s_out<= "10010111";
	WHEN "10000110" => s_out<= "01000100";
	WHEN "10000111" => s_out<= "00010111";
	WHEN "10001000" => s_out<= "11000100";
	WHEN "10001001" => s_out<= "10100111";
	WHEN "10001010" => s_out<= "01111110";
	WHEN "10001011" => s_out<= "00111101";
	WHEN "10001100" => s_out<= "01100100";
	WHEN "10001101" => s_out<= "01011101";
	WHEN "10001110" => s_out<= "00011001";
	WHEN "10001111" => s_out<= "01110011";
	--tenth row
	WHEN "10010000" => s_out<= "01100000";
	WHEN "10010001" => s_out<= "10000001";
	WHEN "10010010" => s_out<= "01001111";
	WHEN "10010011" => s_out<= "11011100";
	WHEN "10010100" => s_out<= "00100010";
	WHEN "10010101" => s_out<= "00101010";
	WHEN "10010110" => s_out<= "10010000";
	WHEN "10010111" => s_out<= "10001000";
	WHEN "10011000" => s_out<= "01000110";
	WHEN "10011001" => s_out<= "11101110";
	WHEN "10011010" => s_out<= "10111000";
	WHEN "10011011" => s_out<= "00010100";
	WHEN "10011100" => s_out<= "11011110";
	WHEN "10011101" => s_out<= "01011110";
	WHEN "10011110" => s_out<= "00001011";
	WHEN "10011111" => s_out<= "11011011";
	--eleventh row	   
	WHEN "10100000" => s_out<= "11100000";
	WHEN "10100001" => s_out<= "00110010";
	WHEN "10100010" => s_out<= "00111010";
	WHEN "10100011" => s_out<= "00001010";
	WHEN "10100100" => s_out<= "01001001";
	WHEN "10100101" => s_out<= "00000110";
	WHEN "10100110" => s_out<= "00100100";
	WHEN "10100111" => s_out<= "01011100";
	WHEN "10101000" => s_out<= "11000010";
	WHEN "10101001" => s_out<= "11010011";
	WHEN "10101010" => s_out<= "10101100";
	WHEN "10101011" => s_out<= "01100010";
	WHEN "10101100" => s_out<= "10010001";
	WHEN "10101101" => s_out<= "10010101";
	WHEN "10101110" => s_out<= "11100100";
	WHEN "10101111" => s_out<= "01111001";
	--twelveth row	    
	WHEN "10110000" => s_out<= "11100111";
	WHEN "10110001" => s_out<= "11001000";
	WHEN "10110010" => s_out<= "00110111";
	WHEN "10110011" => s_out<= "01101101";
	WHEN "10110100" => s_out<= "10001101";
	WHEN "10110101" => s_out<= "11010101";
	WHEN "10110110" => s_out<= "01001110";
	WHEN "10110111" => s_out<= "10101001";
	WHEN "10111000" => s_out<= "01101100";
	WHEN "10111001" => s_out<= "01010110";
	WHEN "10111010" => s_out<= "11110100";
	WHEN "10111011" => s_out<= "11101010";
	WHEN "10111100" => s_out<= "01100101";
	WHEN "10111101" => s_out<= "01111010";
	WHEN "10111110" => s_out<= "10101110";
	WHEN "10111111" => s_out<= "00001000";
	--thirteenth row	    
	WHEN "11000000" => s_out<= "10111010";
	WHEN "11000001" => s_out<= "01111000";
	WHEN "11000010" => s_out<= "00100101";
	WHEN "11000011" => s_out<= "00101110";
	WHEN "11000100" => s_out<= "00011100";
	WHEN "11000101" => s_out<= "10100110";
	WHEN "11000110" => s_out<= "10110100";
	WHEN "11000111" => s_out<= "11000110";
	WHEN "11001000" => s_out<= "11101000";
	WHEN "11001001" => s_out<= "11011101";
	WHEN "11001010" => s_out<= "01110100";
	WHEN "11001011" => s_out<= "00011111";
	WHEN "11001100" => s_out<= "01001011";
	WHEN "11001101" => s_out<= "10111101";
	WHEN "11001110" => s_out<= "10001011";
	WHEN "11001111" => s_out<= "10001010";
	--forteenth row	     
	WHEN "11010000" => s_out<= "01110000";
	WHEN "11010001" => s_out<= "00111110";
	WHEN "11010010" => s_out<= "10110101";
	WHEN "11010011" => s_out<= "01100110";
	WHEN "11010100" => s_out<= "01001000";
	WHEN "11010101" => s_out<= "00000011";
	WHEN "11010110" => s_out<= "11110110";
	WHEN "11010111" => s_out<= "00001110";
	WHEN "11011000" => s_out<= "01100001";
	WHEN "11011001" => s_out<= "00110101";
	WHEN "11011010" => s_out<= "01010111";
	WHEN "11011011" => s_out<= "10111001";
	WHEN "11011100" => s_out<= "10000110";
	WHEN "11011101" => s_out<= "11000001";
	WHEN "11011110" => s_out<= "00011101";
	WHEN "11011111" => s_out<= "10011110";
	--fifteenth row	     
	WHEN "11100000" => s_out<= "11100001";
	WHEN "11100001" => s_out<= "11111000";
	WHEN "11100010" => s_out<= "10011000";
	WHEN "11100011" => s_out<= "00010001";
	WHEN "11100100" => s_out<= "01101001";
	WHEN "11100101" => s_out<= "11011001";
	WHEN "11100110" => s_out<= "10001110";
	WHEN "11100111" => s_out<= "10010100";
	WHEN "11101000" => s_out<= "10011011";
	WHEN "11101001" => s_out<= "00011110";
	WHEN "11101010" => s_out<= "10000111";
	WHEN "11101011" => s_out<= "11101001";
	WHEN "11101100" => s_out<= "11001110";
	WHEN "11101101" => s_out<= "01010101";
	WHEN "11101110" => s_out<= "00101000";
	WHEN "11101111" => s_out<= "11011111";
	--sixteenth row	     
	WHEN "11110000" => s_out<= "10001100";
	WHEN "11110001" => s_out<= "10100001";
	WHEN "11110010" => s_out<= "10001001";
	WHEN "11110011" => s_out<= "00001101";
	WHEN "11110100" => s_out<= "10111111";
	WHEN "11110101" => s_out<= "11100110";
	WHEN "11110110" => s_out<= "01000010";
	WHEN "11110111" => s_out<= "01101000";
	WHEN "11111000" => s_out<= "01000001";
	WHEN "11111001" => s_out<= "10011001";
	WHEN "11111010" => s_out<= "00101101";
	WHEN "11111011" => s_out<= "00001111";
	WHEN "11111100" => s_out<= "10110000";
	WHEN "11111101" => s_out<= "01010100";
	WHEN "11111110" => s_out<= "10111011";
	WHEN "11111111" => s_out<= "00010110";
		     
		     
		     
		     
	WHEN OTHERS => s_out<= "XXXXXXXX";	    
		    
end case;
end process;		    
		    
END beh;			    
			    

